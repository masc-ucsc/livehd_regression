module expression_00181(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(|(|{(~&{(3'd4),(2'd0),(4'sd1)})})),({(5'sd8),(5'sd1),(5'sd12)}!=={{(-2'sd0)}})};
  localparam [4:0] p1 = (((-3'sd1)|(5'd0))===((2'd3)^~(5'sd9)));
  localparam [5:0] p2 = {{4{((3'sd0)!=(3'd7))}}};
  localparam signed [3:0] p3 = (!(^(~^(|(^(((5'd7)===(-2'sd0))^~(+(5'd17))))))));
  localparam signed [4:0] p4 = (^({2{((2'd3)^(5'd1))}}>=(((5'd16)^(4'd15))>>((2'sd0)+(5'd26)))));
  localparam signed [5:0] p5 = ((~&(4'd2 * (^((4'd1)?(2'd1):(3'd0)))))!=(&(((4'sd2)<<(-5'sd2))?((5'd6)?(-2'sd1):(-5'sd12)):((-4'sd2)==(4'd12)))));
  localparam [3:0] p6 = {3{{3{{1{(-2'sd1)}}}}}};
  localparam [4:0] p7 = {(2'd2)};
  localparam [5:0] p8 = (3'sd2);
  localparam signed [3:0] p9 = (+(~|(|(~^(!{2{{3{(-3'sd3)}}}})))));
  localparam signed [4:0] p10 = {3{{3{(3'sd1)}}}};
  localparam signed [5:0] p11 = {({{{(5'sd14)},((4'sd6)?(-3'sd3):(3'd1))}}^~(((5'd6)&&(3'd7))+((3'sd2)>>>(2'd3))))};
  localparam [3:0] p12 = (4'd2 * ((3'd0)<<(3'd3)));
  localparam [4:0] p13 = (-4'sd5);
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = {4{(((-2'sd0)&&(5'd15))<<<((-4'sd0)<=(5'd28)))}};
  localparam signed [4:0] p16 = (+(2'd3));
  localparam signed [5:0] p17 = (+(((-4'sd5)<<(2'd0))+((4'd8)?(5'sd3):(-2'sd0))));

  assign y0 = (((p15^p14)||(!{a1,b1}))<(~^(-4'sd7)));
  assign y1 = ((p13||p5)<<<(p4||b0));
  assign y2 = (-(4'sd1));
  assign y3 = (4'd2 * {4{p14}});
  assign y4 = (a4>b0);
  assign y5 = (((^(a4^~p2))!=(~&(^b0)))|(~(^((p16)>=(+p5)))));
  assign y6 = (((p3!=b0)%p6)<<(((p5==a4)*(p15))));
  assign y7 = {(p4?p2:a4),(5'd9),{4{p8}}};
  assign y8 = (~(-(+(^(4'd7)))));
  assign y9 = (($signed(p3)-(p17>=p8))?((b5^~p14)>>>(-5'sd5)):(p15?a5:p8));
  assign y10 = (5'd2 * (-{1{p13}}));
  assign y11 = (^(^((~^{{a5},(a0>>>a2)})<{(~(b3>>a4))})));
  assign y12 = (~(~&(!((p9?p16:p6)&&(p7?p14:p10)))));
  assign y13 = ((($unsigned(p15)>(4'd13))-(-3'sd2))<<<($signed((-4'sd5))>((a3)>>>(p1+p5))));
  assign y14 = (+{b3,a5,b2});
  assign y15 = (2'd0);
  assign y16 = (|{a3,b5,a4});
  assign y17 = (({{a4,b2},{b2}}+((+a1)&&(-a3)))-(~^(~(~(^{(a3<<b3)})))));
endmodule
