module expression_00363(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{{(3'sd0),(2'd1),(4'd3)}}}==={4{(5'd1)}});
  localparam [4:0] p1 = {(|(-(3'sd1))),(4'd15),((-3'sd1)?(4'sd7):(5'sd11))};
  localparam [5:0] p2 = {2{((5'sd6)!=(3'd1))}};
  localparam signed [3:0] p3 = (((-2'sd1)>=(4'd12))!={4{(5'd17)}});
  localparam signed [4:0] p4 = ({2{((-4'sd6)?(2'd1):(3'd4))}}?(!((5'd3)===(3'sd1))):((2'd3)?(4'd5):(-2'sd0)));
  localparam signed [5:0] p5 = ({1{((4'd5)<<<(5'sd1))}}>=((3'sd0)||(5'd27)));
  localparam [3:0] p6 = (4'd8);
  localparam [4:0] p7 = (&((((5'd15)<<<(4'd5))>(~&(4'sd7)))?(((2'sd0)?(3'sd0):(3'd0))||((-3'sd0)===(3'd7))):(+((-2'sd0)%(-2'sd0)))));
  localparam [5:0] p8 = {4{((5'sd0)-(3'd2))}};
  localparam signed [3:0] p9 = ((-5'sd2)>(-5'sd6));
  localparam signed [4:0] p10 = (|(4'd14));
  localparam signed [5:0] p11 = (2'sd0);
  localparam [3:0] p12 = {2{{4{((-2'sd0)!==(-3'sd0))}}}};
  localparam [4:0] p13 = ((!(+((4'd0)>>>(3'd3))))?(((-2'sd1)>>(4'sd5))>((-3'sd2)<(3'd4))):(((3'sd2)?(-2'sd0):(3'd2))&(|(5'd19))));
  localparam [5:0] p14 = (4'd2 * {((5'd7)>>(4'd15))});
  localparam signed [3:0] p15 = (-4'sd2);
  localparam signed [4:0] p16 = {(((-3'sd1)||(2'd0))<<{1{(3'd0)}}),{4{(4'sd0)}}};
  localparam signed [5:0] p17 = (2'd1);

  assign y0 = {1{((~^(&{1{(^(|p9))}}))?((~&b2)?(~&a3):(|b1)):{3{(^a0)}})}};
  assign y1 = ({(~^a5),{1{b5}},(|b2)}?((b2?b1:p16)?(a0?b5:b2):{p5,p12}):{1{{4{b5}}}});
  assign y2 = (^(((a3<<b5)>>>{b0,b2,b4})>>((b1||a0)>(+a1))));
  assign y3 = ({1{(p12?a1:p5)}}&((2'd3)<<<(p6?p5:b3)));
  assign y4 = (((p16>=p11)-(4'd2 * a0))<<<((&(p11|p11))!=(b3===b2)));
  assign y5 = (5'd15);
  assign y6 = ({2{(~&(p14>=p11))}}<<({4{p11}}?(p6?b5:p4):{2{p6}}));
  assign y7 = ((|p1)^~(p14-p10));
  assign y8 = {4{(3'd5)}};
  assign y9 = {2{(3'd0)}};
  assign y10 = (((^(^p12))?(|(|p11)):{3{p6}})<(|{(^(-{2{p10}})),({p6,p0,p12}<=(a3!=p2))}));
  assign y11 = (6'd2 * $unsigned(p10));
  assign y12 = $unsigned({(p4+b2)});
  assign y13 = (+((^(-4'sd7))%a0));
  assign y14 = (a4<<<p7);
  assign y15 = (!{4{(|(-5'sd15))}});
  assign y16 = (5'd19);
  assign y17 = (((p2-p2))<((p15)^(4'sd1)));
endmodule
