module expression_00928(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(4'sd7));
  localparam [4:0] p1 = {1{((5'd11)?(3'sd0):(-4'sd4))}};
  localparam [5:0] p2 = (2'd3);
  localparam signed [3:0] p3 = ((4'sd2)&(5'd23));
  localparam signed [4:0] p4 = {3{(((-5'sd12)^(2'sd1))&(-2'sd0))}};
  localparam signed [5:0] p5 = (4'd14);
  localparam [3:0] p6 = {3{((4'd13)-(-2'sd0))}};
  localparam [4:0] p7 = ({1{({2{(3'd5)}}!=((5'd23)?(-4'sd6):(-4'sd3)))}}>>{{(-4'sd3),(2'd1)},((3'sd1)?(4'sd1):(4'sd7))});
  localparam [5:0] p8 = ((5'd25)?(5'sd15):(-2'sd1));
  localparam signed [3:0] p9 = ((5'd31)^~(-5'sd5));
  localparam signed [4:0] p10 = (((5'd16)+(|(3'sd0)))===(3'sd1));
  localparam signed [5:0] p11 = ((((3'd5)?(4'd14):(5'd24))?{(3'sd2),(-5'sd11)}:((-4'sd3)<(3'sd3)))!=({(-2'sd0),(4'd15)}?((4'sd0)?(2'sd1):(3'd1)):{(3'sd3),(3'd1),(2'sd1)}));
  localparam [3:0] p12 = (-(~|(-4'sd7)));
  localparam [4:0] p13 = ((((4'sd3)?(4'd0):(4'd10))<<((~(5'sd14))>>((2'd3)<(3'd2))))<<(((4'sd2)!==(5'd23))?(^((3'd5)?(-5'sd1):(3'sd1))):((5'd27)<=(5'd12))));
  localparam [5:0] p14 = (((2'd2)?(-3'sd0):(3'sd2))>=((^(4'd9))&((5'd21)?(3'd0):(3'd4))));
  localparam signed [3:0] p15 = ((2'sd1)>(3'sd3));
  localparam signed [4:0] p16 = (((4'd2)?(2'sd1):(5'sd11))?((-5'sd8)?(4'sd6):(-3'sd0)):((3'd7)?(5'd11):(4'd9)));
  localparam signed [5:0] p17 = (-5'sd15);

  assign y0 = (((-4'sd4))+((5'd2 * $unsigned((p2^~a2)))<{2{(p10)}}));
  assign y1 = (4'sd5);
  assign y2 = (2'd2);
  assign y3 = (|{4{{1{(~|a5)}}}});
  assign y4 = ({(2'sd0)});
  assign y5 = ((p11<=a3)>(a0));
  assign y6 = (({a1,p4,b4}>>>(^{b4,b3}))<=(+({b4,b1}>>>(~a1))));
  assign y7 = (b2|b1);
  assign y8 = {(p17>p16),(p8?p5:p0),{p7,p17,p5}};
  assign y9 = (p7>p13);
  assign y10 = ((~&p10)||(&b4));
  assign y11 = ((({p15,b5,p2}|{p1})>>>({p5}||(p1>>p6)))>{((5'd17)||((4'sd5)>>>{b3}))});
  assign y12 = (((p1%p13)%a1)+((b1!==b0)<<<(p6<=p5)));
  assign y13 = (({a2,a1,b0}&&(-5'sd2))?{(~&a1),(a5<p8),$signed(p10)}:((|a2)?(5'd0):(p2?b3:a4)));
  assign y14 = (p17?p1:p12);
  assign y15 = ((p1?p17:p6)?$signed(p2):(p16&&p13));
  assign y16 = (-5'sd0);
  assign y17 = {(a1<=a4),{(b3-a2)}};
endmodule
