module expression_00259(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd13);
  localparam [4:0] p1 = (~(5'd27));
  localparam [5:0] p2 = ((((5'd31)?(5'd16):(4'd13))<={(2'd1),(2'sd1)})!==(((-4'sd3)&(2'sd0))>>>(~(3'd2))));
  localparam signed [3:0] p3 = (3'd4);
  localparam signed [4:0] p4 = {3{(3'd0)}};
  localparam signed [5:0] p5 = (^(~|((2'sd0)===(4'd3))));
  localparam [3:0] p6 = (({((-2'sd1)?(3'd1):(3'd6)),((2'd3)?(3'sd1):(2'd2))}<<<(4'd12))>={({(3'd6),(2'd3)}?((4'sd4)?(3'd5):(4'sd1)):((4'd3)?(3'sd0):(-5'sd1)))});
  localparam [4:0] p7 = ((~|(((3'sd2)!==(4'd5))>{(2'd0)}))?(((-3'sd2)<<<(-2'sd1))||((3'sd1)==(3'd0))):(~^{4{(5'd29)}}));
  localparam [5:0] p8 = ((6'd2 * (5'd23))<<(~&(5'sd4)));
  localparam signed [3:0] p9 = (((-2'sd0)>=(5'd17))?((4'd3)&&(-3'sd1)):{2{(2'd2)}});
  localparam signed [4:0] p10 = {(5'd28),(4'd7),(-2'sd0)};
  localparam signed [5:0] p11 = ((~&({(2'd1),(-5'sd2)}+(&(3'sd1))))&((~^(5'sd5))>=(^(3'd0))));
  localparam [3:0] p12 = (((-2'sd0)?(4'd4):(3'd4))?((-2'sd1)?(5'd11):(4'd11)):((4'd11)-(-5'sd8)));
  localparam [4:0] p13 = {({2{(5'd12)}}?((2'sd0)?(-3'sd0):(4'sd6)):((5'd14)?(5'd26):(-5'sd4))),(((-2'sd0)?(2'd0):(5'd28))?{2{(2'd3)}}:{(-2'sd1)}),{3{((3'd4)?(-3'sd3):(5'd22))}}};
  localparam [5:0] p14 = ({1{{1{(^(4'd3))}}}}?(!(-4'sd6)):(((5'sd6)-(3'd4))+{(5'd29),(-5'sd9)}));
  localparam signed [3:0] p15 = (~^((6'd2 * (-(+(3'd3))))>>(((2'd0)&&(5'sd8))!=((-4'sd0)&(-4'sd6)))));
  localparam signed [4:0] p16 = ((4'sd2)?(5'sd4):((2'sd1)?(-2'sd0):(5'sd4)));
  localparam signed [5:0] p17 = ((((-2'sd1)==(-4'sd6))^~((-2'sd1)+(5'd13)))>>>(!(((2'd0)/(4'sd3))/(2'd3))));

  assign y0 = (((b4?a1:b2)?{p7,b0}:{a1,b1})<(((p8!=a4)==(a0))==((b4&a0)||(a4<<p6))));
  assign y1 = ((-b2)?(a2^a1):(~|p5));
  assign y2 = (4'sd3);
  assign y3 = (2'sd1);
  assign y4 = (~&(((b4|p10)?(3'sd3):(|b5))<<<(!(2'sd1))));
  assign y5 = (&(+((-(-3'sd3))!==(b3>>>b0))));
  assign y6 = {3{(!(~&(&p1)))}};
  assign y7 = (({(p2^a3)}>(2'sd1))>>>{(3'd4),(5'd31),(3'd6)});
  assign y8 = {2{b3}};
  assign y9 = ((p1?p1:b4)>>(p8?a5:a1));
  assign y10 = {4{(3'sd1)}};
  assign y11 = $unsigned((^{3{{(~^(|a0)),({3{a1}})}}}));
  assign y12 = $signed((-5'sd2));
  assign y13 = (^(({b4,b5}<<<$unsigned({b3,a1}))<=(|(~{{b5},{a5,a3}}))));
  assign y14 = (((2'sd1)>>>(4'd2 * (b1&&a1)))===(~|(5'sd2)));
  assign y15 = (a2>=b1);
  assign y16 = $unsigned((((a3+a2)===(&b4))?{(a2>>a2),(a0?a3:b1)}:({p16,a3,b0}>=(a2>>b2))));
  assign y17 = {(a3?p12:b0),{2{a5}}};
endmodule
