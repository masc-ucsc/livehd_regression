module expression_00762(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd1);
  localparam [4:0] p1 = (((2'sd1)?(4'sd3):(4'd12))!=(((5'd12)?(5'sd8):(5'sd0))*((4'd9)?(-5'sd0):(5'd21))));
  localparam [5:0] p2 = (((2'd1)+(-3'sd1))>>(~((-4'sd7)&&(-5'sd10))));
  localparam signed [3:0] p3 = ((5'd1)<<(-3'sd3));
  localparam signed [4:0] p4 = ((|(-2'sd0))^~((3'd2)^~(4'sd0)));
  localparam signed [5:0] p5 = (^{(((4'd12)<(5'sd3))<(~(2'sd1)))});
  localparam [3:0] p6 = ((!(5'd2 * {4{(2'd1)}}))&(~&(-(3'sd0))));
  localparam [4:0] p7 = (((+(3'sd3))<<(^(4'd0)))!=(4'd9));
  localparam [5:0] p8 = {2{(!{2{{(3'd7),(4'd8)}}})}};
  localparam signed [3:0] p9 = (+(~|(~|((~(~&(-4'sd0)))+(~|(+(3'sd1)))))));
  localparam signed [4:0] p10 = (|((3'sd0)>>(-4'sd6)));
  localparam signed [5:0] p11 = {4{{1{(-4'sd2)}}}};
  localparam [3:0] p12 = ((|(~(-5'sd14)))^((3'd4)===(5'sd15)));
  localparam [4:0] p13 = {((((2'sd0)!=(3'd5))<(~&(4'sd7)))^~(~^(((-4'sd1)>(3'd4))||{1{(5'd11)}})))};
  localparam [5:0] p14 = {{((2'sd1)?(2'd3):(2'd1))}};
  localparam signed [3:0] p15 = ({{{{(-2'sd0),(3'd5),(3'sd1)},((-5'sd2)-(-2'sd1)),((3'd2)-(2'sd0))}}}<<{{4{{3{(-3'sd2)}}}}});
  localparam signed [4:0] p16 = (((4'sd3)?(3'd0):(-4'sd6))?(((-3'sd0)?(5'sd6):(-5'sd14))!=(^(3'd2))):(5'sd9));
  localparam signed [5:0] p17 = (3'd2);

  assign y0 = $unsigned((~^p17));
  assign y1 = ((((a5^b4)|{a1}))-{($signed({p10,b4}))});
  assign y2 = $unsigned((3'd6));
  assign y3 = ((b0/a5)>>>(b1/a2));
  assign y4 = (^(!(~&({((~|(+a1))<<(b2^~b2))}^~((b4==a0)^(-{b4,b4}))))));
  assign y5 = {4{{4{b0}}}};
  assign y6 = (((a1?b3:b0)===({3{a5}}<(a5&a2)))&&((!(p14>p0))?(b5!==a1):(p14<=p2)));
  assign y7 = (-5'sd7);
  assign y8 = {(2'd2),(&(-((b2?a1:p9)<<<{p3,p13,p12})))};
  assign y9 = (((p15!=b4)?(p3*p8):(p5>>>p6))<<<((p11?p6:p16)?(p17?b4:p17):(~&p1)));
  assign y10 = {b5,p14,p4};
  assign y11 = {4{{4{a2}}}};
  assign y12 = (~&{1{a0}});
  assign y13 = {p4,p11,b1};
  assign y14 = {(-({1{(-(&(~|(~|{p12,a5,p10}))))}}))};
  assign y15 = (~&p10);
  assign y16 = (4'd7);
  assign y17 = {3{(4'sd0)}};
endmodule
