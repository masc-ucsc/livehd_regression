module expression_00852(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{({((3'd4)?(2'sd1):(4'd12))}?(!(~|((4'd14)|(3'd5)))):((5'sd13)?(3'sd2):(5'd17)))}};
  localparam [4:0] p1 = (2'd2);
  localparam [5:0] p2 = ((-3'sd2)/(5'd17));
  localparam signed [3:0] p3 = (((5'd12)===(5'd11))^((2'd0)>=(2'd2)));
  localparam signed [4:0] p4 = (((2'd1)?(2'd1):(-2'sd0))?(5'd2 * (2'd0)):{{(-5'sd2)}});
  localparam signed [5:0] p5 = ((!(((5'sd2)?(2'd0):(5'd16))||((2'd0)<(3'd6))))^(-(!((-3'sd1)?(2'sd1):(3'd0)))));
  localparam [3:0] p6 = (&(4'd6));
  localparam [4:0] p7 = (^(-((|{3{(5'sd8)}})<{(4'd10),(4'sd3),(-3'sd3)})));
  localparam [5:0] p8 = (~^(|(5'd11)));
  localparam signed [3:0] p9 = (4'd4);
  localparam signed [4:0] p10 = ((3'sd1)<<(2'd1));
  localparam signed [5:0] p11 = {(({(3'd0),(4'd12)}>>>{(2'd3)})>=(-{((-3'sd1)>>(-2'sd0)),((-2'sd0)>(-2'sd0))}))};
  localparam [3:0] p12 = (&((~&(3'd0))!==((-2'sd1)<<(-5'sd9))));
  localparam [4:0] p13 = {{((2'd0)&&(-3'sd1)),{(3'd5),(4'd10),(3'd1)}}};
  localparam [5:0] p14 = (((2'd2)>>(4'd1))!=={1{(4'sd3)}});
  localparam signed [3:0] p15 = (&{2{{4{((-2'sd0)-(5'd13))}}}});
  localparam signed [4:0] p16 = ((-5'sd8)<(3'd6));
  localparam signed [5:0] p17 = (|(+{2{{4{(~^(4'd4))}}}}));

  assign y0 = (3'sd0);
  assign y1 = (+(5'd2 * (4'd3)));
  assign y2 = ((~&(5'sd1))<(+((-(~&{b4,b5,p1}))&&((-3'sd3)+(3'd1)))));
  assign y3 = {3{(~&(b0?a0:a3))}};
  assign y4 = (a5^p9);
  assign y5 = {((5'd2 * $unsigned(p5)))};
  assign y6 = (((a1||a3)|(b0==p5))?((a0&&a5)&&(a3|b4)):{1{(b1|p5)}});
  assign y7 = (~&{$unsigned($unsigned((~^$signed({b4,b4,a1})))),$unsigned($signed({(5'd16),(a5),{b1,a0}}))});
  assign y8 = ((!{(a3>>a4),(b5?b2:b4),(a1>>>a2)})!==(2'sd1));
  assign y9 = (-2'sd1);
  assign y10 = ($unsigned((p8>=p15))?$signed((p13?p1:p7)):(2'd0));
  assign y11 = ((5'd5)<<<(5'sd6));
  assign y12 = {3{{p3,p6,p6}}};
  assign y13 = {4{(p0?p9:p17)}};
  assign y14 = $signed((~(~(((p2<p10)*(a1?p6:a0))?(~(~^(b4>=p13))):(b5?p1:p10)))));
  assign y15 = (-((&((a5/b1)>>>(a0||a0)))|(!(((p2>b5)^((4'd0)))))));
  assign y16 = {{{{p10,p12,b5},{b4},{b0}}},{{{p4,a0},{b2,b0}}},{{b0,b0},{b5,a3,p12}}};
  assign y17 = (((-b3)<<(a2>=a3))!==(~(&{b0,b1})));
endmodule
