module expression_00538(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~((4'sd5)<=(4'd10)));
  localparam [4:0] p1 = (~|{{(3'd7),(5'sd12)}});
  localparam [5:0] p2 = (((4'd13)?(2'd2):(2'd1))?(4'd5):((5'd2 * (2'd2))<=((5'sd10)<=(4'd6))));
  localparam signed [3:0] p3 = {(4'sd1),(5'd1)};
  localparam signed [4:0] p4 = {(^(^(4'd11))),{2{(-3'sd0)}}};
  localparam signed [5:0] p5 = (~&{2{{2{(3'd4)}}}});
  localparam [3:0] p6 = (!{{(-2'sd1),(3'd4),(5'sd14)},(-(3'd1)),{(3'd5),(3'd2)}});
  localparam [4:0] p7 = {(2'd0),(2'sd1),(4'd8)};
  localparam [5:0] p8 = ({4{(5'sd10)}}<(-4'sd3));
  localparam signed [3:0] p9 = (((-2'sd0)>(4'sd4))%(4'd14));
  localparam signed [4:0] p10 = ({2{((-5'sd11)&&(-3'sd0))}}||({1{(5'd16)}}>>>((4'sd5)==(-4'sd4))));
  localparam signed [5:0] p11 = ((&((-5'sd7)?(4'sd5):(2'sd1)))?(^(~^(-4'sd6))):((4'sd6)>>(2'd2)));
  localparam [3:0] p12 = ({((5'd2 * (2'd1))<=((-5'sd13)?(-3'sd2):(2'd0)))}<<<{{(4'sd2),(3'sd2)},((-5'sd4)?(-4'sd5):(4'sd3)),((2'd0)^(-4'sd2))});
  localparam [4:0] p13 = ((3'd0)?(4'd1):(4'sd5));
  localparam [5:0] p14 = (~&(((3'sd3)&((-3'sd0)<(5'd17)))&&(-(3'd4))));
  localparam signed [3:0] p15 = ((2'd3)?(-4'sd1):(-3'sd1));
  localparam signed [4:0] p16 = {2{((-3'sd0)?(4'd3):(-4'sd1))}};
  localparam signed [5:0] p17 = (((-2'sd0)?(5'd22):(-3'sd1))?({1{(5'sd2)}}!=((3'sd0)&&(4'd14))):({2{(5'd31)}}^~((3'd1)?(-2'sd1):(-5'sd5))));

  assign y0 = (~&((-(^(|(((&(a2?p17:a4))?(~&(~^b3)):(~^$signed(a3)))))))));
  assign y1 = $unsigned({((p0?p6:b3)^{p10,p10}),{(p17),(5'sd12),{a2}},({p7,p17}+(p10^p5))});
  assign y2 = (~|((~(|a1))/a0));
  assign y3 = ((p7>>p15)!=(^(p0&&p17)));
  assign y4 = ((-3'sd2)>=(~({(5'd11)}>((3'd3)^(5'd9)))));
  assign y5 = ((p9>>>p8)*(2'sd1));
  assign y6 = (3'd5);
  assign y7 = ((~(&((!((~|b1)<(~^a1))))))<<(($unsigned(p1)<<(!b5))^~(^(p1<=a1))));
  assign y8 = {{(4'd2 * {1{{p1}}}),((p10?p2:p17)-(p16?p9:p8))}};
  assign y9 = (~&(-$signed($unsigned($unsigned(((((+(~|$unsigned($signed(b5))))))^((((~|a5))!==$signed((~|a3))))))))));
  assign y10 = (~&(!{4{{{2{a2}},(!b4),{b1,p11,b3}}}}));
  assign y11 = (3'd7);
  assign y12 = {(p6^~a1)};
  assign y13 = (+{2{((p11-p14)>=(-2'sd0))}});
  assign y14 = ((((4'sd6)<=(-3'sd0))>>>(-4'sd4))+(5'sd7));
  assign y15 = (-4'sd2);
  assign y16 = (((a4&p9)-(6'd2 * p8))?((b4<<<p9)!=(p10>>>p11)):((p15>>p1)<=(p8?p17:b0)));
  assign y17 = (2'sd1);
endmodule
