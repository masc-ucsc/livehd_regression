module expression_00942(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{{3{((-2'sd1)<=(2'd0))}}}};
  localparam [4:0] p1 = ((-3'sd2)&&(3'd3));
  localparam [5:0] p2 = (-2'sd1);
  localparam signed [3:0] p3 = ((-5'sd0)>>>({1{{3{(4'd9)}}}}^{2{(3'd4)}}));
  localparam signed [4:0] p4 = ({{(4'sd1),(3'd3)},((-5'sd7)<<<(-3'sd3)),((5'sd6)>>>(-4'sd2))}===({(5'd21),(5'd29),(2'd2)}>>{(4'sd2),(5'sd8),(2'sd0)}));
  localparam signed [5:0] p5 = {1{(~|(5'd18))}};
  localparam [3:0] p6 = {1{(4'd13)}};
  localparam [4:0] p7 = ((|((|(4'd8))&(5'd2 * (2'd0))))&&(((-5'sd14)&(2'd0))+{3{(4'd6)}}));
  localparam [5:0] p8 = ((~((-5'sd3)?(5'd19):(4'd15)))?(((-3'sd3)>(3'd6))&&((3'd2)?(5'd14):(4'sd1))):{{4{(4'sd6)}},(+(-4'sd7)),(3'sd1)});
  localparam signed [3:0] p9 = (~|(((-4'sd3)?(3'd6):{(5'd30),(-2'sd0),(-2'sd1)})===((4'sd1)<<<(5'sd9))));
  localparam signed [4:0] p10 = (2'sd1);
  localparam signed [5:0] p11 = {4{{4{(-2'sd1)}}}};
  localparam [3:0] p12 = {{2{{{((4'sd5)^(-4'sd2)),((-4'sd6)!=(-4'sd3))}}}}};
  localparam [4:0] p13 = ((5'd13)?(-{4{(-2'sd1)}}):(-5'sd0));
  localparam [5:0] p14 = {3{(5'd4)}};
  localparam signed [3:0] p15 = (~^(~&(-((((4'sd3)===(-5'sd9))|((5'd18)&(-5'sd8)))<(^((3'd6)+(5'd4)))))));
  localparam signed [4:0] p16 = (+((|(|((|(2'd2))^~((2'd2)>>(2'd1)))))>=((!(~^(5'd16)))|(~(~&(5'd29))))));
  localparam signed [5:0] p17 = {((((4'd12)?(2'd2):(2'd2))&{(5'd27)})&&(((5'd10)<=(2'sd1))>{(-4'sd5),(-4'sd5),(-5'sd2)}))};

  assign y0 = {a3,b5};
  assign y1 = ((~|$unsigned({b5,a2}))===((b0-b2)!=(~a2)));
  assign y2 = (4'sd0);
  assign y3 = ((|b2)?(p6?p9:p17):(5'd11));
  assign y4 = {2{((a5?b0:b1)^(p5?b4:p12))}};
  assign y5 = (&(6'd2 * (b1>=p6)));
  assign y6 = (6'd2 * (a1/a0));
  assign y7 = (^(((a3!==a0)?(~|{p10,a0,p2}):{a0,b2})^({b4,a4}?(!(b3-p16)):(a4?b0:p12))));
  assign y8 = (~^(~^((~^((^b4)&(p1?p3:b0)))>>>(~&(6'd2 * (~(|a2)))))));
  assign y9 = ((5'sd13)!=((p3>>>p14)^~(p13/b5)));
  assign y10 = (~(|(+((4'd11)&((+(p15>>p13))<<(&(4'd4)))))));
  assign y11 = (~|$signed((~&$unsigned($signed((~&(-(!($signed((((((|((~^a0)))))))))))))))));
  assign y12 = (({{b5,a0},(+p16)}>>>((p3&&p6)<<{p11}))||({4{a1}}!={{4{p15}},{b1,p1,p3}}));
  assign y13 = {{3{p5}},(p10?p9:p2)};
  assign y14 = ({1{$signed(((a1?b3:b1)?{2{b2}}:$unsigned((a0?b5:b5))))}}==({2{a4}}?(a3?a1:a2):((b4?b3:b0))));
  assign y15 = $unsigned((~|{4{{1{(-(a1))}}}}));
  assign y16 = {4{((p5<<<p12))}};
  assign y17 = ((b3==a3)?(4'sd1):(b3?a4:b5));
endmodule
