module expression_00817(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{({2{(5'd2)}}+{4{(5'sd0)}})},(((4'd13)>(4'd8))>>>((5'd15)!==(2'd1)))};
  localparam [4:0] p1 = (!(^{{(3'sd1),(5'd18)}}));
  localparam [5:0] p2 = {{(2'd2),(2'd1),(2'd1)},((5'sd10)<<(5'sd12)),(-((3'd4)?(-3'sd3):(-3'sd2)))};
  localparam signed [3:0] p3 = ((5'd2 * (^(2'd1)))?(^((3'd2)+(3'd1))):((4'd7)?(3'd7):(2'd1)));
  localparam signed [4:0] p4 = (-(5'sd15));
  localparam signed [5:0] p5 = {1{(+{1{(~&(~(&(~|(4'd3)))))}})}};
  localparam [3:0] p6 = (~^(~^({4{{2{(3'd4)}}}}|((~(-4'sd3))?{(4'd9),(4'd4),(4'd4)}:((3'd3)>=(-2'sd0))))));
  localparam [4:0] p7 = (-{2{({4{(4'd0)}}>>>(-((2'd3)-(3'd1))))}});
  localparam [5:0] p8 = (5'd22);
  localparam signed [3:0] p9 = (^(3'd1));
  localparam signed [4:0] p10 = ((-2'sd1)-(5'd7));
  localparam signed [5:0] p11 = ((-4'sd0)==(4'd6));
  localparam [3:0] p12 = ({(((4'd5)&(3'sd1))<<(-{(2'd0),(2'd3),(-3'sd0)}))}<<((&((-2'sd0)<<(4'sd4)))>>>(~&(~|(5'sd0)))));
  localparam [4:0] p13 = ((3'd2)?(5'sd7):(5'd22));
  localparam [5:0] p14 = ({(5'd24),(3'd1),(2'd0)}?{(3'sd0)}:((2'sd0)?(3'd1):(2'd3)));
  localparam signed [3:0] p15 = {((4'd4)>=((-5'sd15)<<(4'sd5))),((!(~|(4'd11)))>(-2'sd0))};
  localparam signed [4:0] p16 = ((&(!(~(2'd3))))>>(|(|(|(3'sd2)))));
  localparam signed [5:0] p17 = ({3{((-5'sd0)!=(5'sd10))}}==(5'd23));

  assign y0 = (~$signed(({2{({4{b2}}>(a1^~b1))}}>>>((!(b1===a0))!=(-(a1+p4))))));
  assign y1 = (|(((b5!==b4)===(b5>>>b0))>>((a5>>>b4)/a5)));
  assign y2 = (+(|(~&(-3'sd3))));
  assign y3 = {3{p11}};
  assign y4 = ({1{(^(3'sd1))}}?((a1?p2:p17)<<<(a0?a3:p8)):(b3?a0:b5));
  assign y5 = {((p10?p1:p11)>>>(p9?p13:p7)),((2'sd0)),(~({p3,p17,p6}<<<(5'd22)))};
  assign y6 = ({3{{2{p6}}}}+(^(~(((5'd13)^{3{b4}})^((b2<<<p11)==(p12<p12))))));
  assign y7 = ((b5?p5:p13)-(p6<<p12));
  assign y8 = {1{{1{(((&p5)>(b1&b0))>=(+(~&(|(p1&p15)))))}}}};
  assign y9 = ((((6'd2 * p14))?(2'd3):(b1!==b3))-((4'd8)!==((3'd6)?(b2===b5):(b1?a4:a4))));
  assign y10 = (5'd23);
  assign y11 = ({3{((p7?p2:p13))}}&&{3{(-{p5,p10,p4})}});
  assign y12 = ({2{{4{p14}}}}>>>({2{p8}}?{p5,p0,p15}:{p13,b1,p2}));
  assign y13 = ((({4{b3}}>>>{2{a4}})^~({1{a2}}^(b1>>a1)))&(({3{b4}}^{4{a4}})<<((p9>>a0)^~{1{b2}})));
  assign y14 = ($signed(p13)&(p7^a4));
  assign y15 = {1{((3'sd2)<<<{2{{3{p7}}}})}};
  assign y16 = (~^((b2?a1:b1)?{(^b4),$signed(b0)}:{(&$unsigned(b1))}));
  assign y17 = (((b0+p0)?(p9):(p6?p2:p5))?((p8?p16:b3)?(b4===b2):$unsigned(p1)):({p10,p11}?{a3}:$signed(p13)));
endmodule
