module expression_00390(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(^((5'd22)?(-5'sd12):(5'sd9))),(|(!(|(2'sd1))))};
  localparam [4:0] p1 = {4{((2'd3)&(-5'sd9))}};
  localparam [5:0] p2 = {4{((2'd1)?(4'd11):(3'd4))}};
  localparam signed [3:0] p3 = (|(4'd6));
  localparam signed [4:0] p4 = (~^(~&(-((3'd1)==(3'd5)))));
  localparam signed [5:0] p5 = (+(4'sd2));
  localparam [3:0] p6 = (((~&(4'sd1))!=={1{(4'd9)}})&(4'sd5));
  localparam [4:0] p7 = (-(~&(5'd17)));
  localparam [5:0] p8 = ((-3'sd1)&&((^((3'd7)-(5'sd0)))<<<((3'd0)>(5'sd5))));
  localparam signed [3:0] p9 = ((5'd2 * (-(5'd20)))!=(((3'd6)?(2'd1):(5'sd0))!=((-5'sd0)?(4'd13):(-3'sd0))));
  localparam signed [4:0] p10 = ((~&(2'd2))&(&(5'd26)));
  localparam signed [5:0] p11 = ({((-4'sd3)-(5'd31)),(~^(3'sd3))}&{(2'd0),(3'sd1),(-4'sd5)});
  localparam [3:0] p12 = (5'd2 * {3{(3'd0)}});
  localparam [4:0] p13 = (~(^(|(|({4{(2'd0)}}&&{1{(5'd2 * ((2'd0)<(4'd9)))}})))));
  localparam [5:0] p14 = ((-4'sd0)?(3'sd3):(4'd11));
  localparam signed [3:0] p15 = (~&(-(^{3{(~(-3'sd3))}})));
  localparam signed [4:0] p16 = (-((!((3'd5)>>(5'd19)))%(5'sd6)));
  localparam signed [5:0] p17 = ({2{{(~(5'd7))}}}>>{((-2'sd0)&&(|(-4'sd5)))});

  assign y0 = {((~^{a2,b0})>>>(4'd8)),(4'd2)};
  assign y1 = $signed(({({p0,p1,p16}&&(2'sd0)),$signed({2{({p5,p1,a4})}})}));
  assign y2 = {p13,p9,p15};
  assign y3 = (((b2>b4)?(a1!=a2):(a3?p0:a0))?{4{(b4?p14:b2)}}:({2{p5}}+$unsigned((b0^~a3))));
  assign y4 = (((2'd1)>=(^(p17)))|((~&(b3?p15:a4))+$signed((a4!==b1))));
  assign y5 = (+(((^(5'd25)))));
  assign y6 = {(3'sd2),(!((a0>=a1)<<<(5'd0))),((2'd2)>>>(-2'sd1))};
  assign y7 = {3{(~|a5)}};
  assign y8 = {2{(-3'sd0)}};
  assign y9 = (!$unsigned($signed($signed($unsigned((&(~^{2{{2{(p2)}}}})))))));
  assign y10 = ((a5<b1)<<{1{b0}});
  assign y11 = {3{b2}};
  assign y12 = (^($signed((p16?b1:p6))<<(!(p12>=p4))));
  assign y13 = {(($signed((((-5'sd2)<<<(-5'sd1))>>>{(p9&&a4),(a4)}))&&(((b1>=a1)>>>(a0&a5))^~(4'd10))))};
  assign y14 = {4{$unsigned(p16)}};
  assign y15 = (4'd0);
  assign y16 = (b1?a3:a2);
  assign y17 = (5'sd0);
endmodule
