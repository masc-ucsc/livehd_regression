module expression_00475(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd1),(-5'sd4)};
  localparam [4:0] p1 = (4'd8);
  localparam [5:0] p2 = ({{(4'd4),(4'd4),(4'sd4)},(2'd3)}>>>(4'd5));
  localparam signed [3:0] p3 = ((~|(((4'd7)||(4'd3))|{1{(4'd13)}}))?({4{(-5'sd1)}}?((5'd17)?(3'd6):(3'sd2)):{(-2'sd0),(3'd6),(5'd14)}):{3{((-5'sd4)>(3'sd3))}});
  localparam signed [4:0] p4 = ((-5'sd2)?(-4'sd4):(3'd5));
  localparam signed [5:0] p5 = (~&({1{{((4'd11)?(3'sd2):(-4'sd5)),{(5'd20)}}}}^{(+((4'd14)||(2'sd1)))}));
  localparam [3:0] p6 = (5'd2 * ((5'd14)^~(2'd0)));
  localparam [4:0] p7 = (&(2'd3));
  localparam [5:0] p8 = (((2'd0)?(2'd2):(5'd16))<<({4{(3'sd3)}}<<((2'sd0)>>(-4'sd4))));
  localparam signed [3:0] p9 = {1{(((3'sd3)>=(4'd2 * (5'd15)))<(4'sd5))}};
  localparam signed [4:0] p10 = (((5'sd11)>(4'd13))^(3'd0));
  localparam signed [5:0] p11 = (~|(4'd2));
  localparam [3:0] p12 = ({(~|(3'sd1))}>>>((2'd2)<=(-3'sd2)));
  localparam [4:0] p13 = {(6'd2 * (3'd7)),{(2'd0),(3'd2)},((-3'sd0)!==(-2'sd1))};
  localparam [5:0] p14 = {3{{4{(-3'sd0)}}}};
  localparam signed [3:0] p15 = ((((3'd1)<<<(2'd2))!=((4'd8)?(2'sd1):(4'sd0)))!=(((4'd10)<=(-4'sd6))>>>((-3'sd1)?(-5'sd6):(3'd2))));
  localparam signed [4:0] p16 = ((~|(|(|(|(2'd3)))))?(^((2'd3)||((4'd12)/(3'd7)))):(!((2'd3)?(-4'sd2):(4'd7))));
  localparam signed [5:0] p17 = (|(-3'sd2));

  assign y0 = ((~^(&((b1||p5)&{4{p6}})))||(~|({4{p15}}^~(p0|p14))));
  assign y1 = {$signed((~(p12?p17:p1))),{3{p16}},((p8?p0:a1))};
  assign y2 = {1{(-{2{(~(~&((^(~p12))^~{1{$unsigned(a3)}})))}})}};
  assign y3 = $signed({{(~|((a4)>>(|p7))),((^b2)>>(~a0)),{{1{a4}},(p6&p4)}}});
  assign y4 = (|(((p14!=p9)-(p15|p17))<=((p15&&p4)<=(p7+b3))));
  assign y5 = (p6^~p13);
  assign y6 = (5'd2 * (~^{1{b1}}));
  assign y7 = ($signed(($unsigned(p0)-(p15!=p0)))>>>($unsigned((b3))>>>((p1||p6))));
  assign y8 = (((!p14)?(a3&&a0):{a1})<<((b4&&p10)?(a0<b2):(a5>>a2)));
  assign y9 = {({p7,p11}|(b2>>>p3)),((p8+p14)<<<{p15}),(a0?a1:p6)};
  assign y10 = ((2'd0)?{{3{b1}}}:(b1?b1:p4));
  assign y11 = (((b5-a2)>>>(b2?b0:a1))>>(-4'sd6));
  assign y12 = (5'd13);
  assign y13 = (4'd14);
  assign y14 = ({3{b0}}<=(a1?b3:b3));
  assign y15 = (~^(2'd0));
  assign y16 = (&((~&((|b5)||{3{p1}}))>>{3{(b5<p6)}}));
  assign y17 = (!(2'd0));
endmodule
