module expression_00060(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd3)<<(4'sd0))%(4'd7))||(((4'd4)===(-4'sd3))!=((2'sd1)^~(5'd21))));
  localparam [4:0] p1 = (4'd3);
  localparam [5:0] p2 = ((|((3'd5)?(3'd1):(3'd4)))===(|((4'd3)==(4'd14))));
  localparam signed [3:0] p3 = (-2'sd1);
  localparam signed [4:0] p4 = (~|((5'd1)?(-5'sd10):(3'sd0)));
  localparam signed [5:0] p5 = {3{((-2'sd1)<<(5'd22))}};
  localparam [3:0] p6 = ((^((3'd2)?(-2'sd1):(2'sd0)))?((2'd3)?(3'sd2):(-5'sd7)):((3'd5)?(4'd14):(-4'sd5)));
  localparam [4:0] p7 = (^((5'sd2)?(5'd21):(-5'sd2)));
  localparam [5:0] p8 = (4'd1);
  localparam signed [3:0] p9 = (3'sd1);
  localparam signed [4:0] p10 = (|(-(-4'sd7)));
  localparam signed [5:0] p11 = {2{{3{{2{(-2'sd0)}}}}}};
  localparam [3:0] p12 = ({3{((-4'sd6)!=(4'd11))}}>=(5'd17));
  localparam [4:0] p13 = {3{(-4'sd7)}};
  localparam [5:0] p14 = ((-(-4'sd2))^((4'd11)?(5'sd5):(-2'sd1)));
  localparam signed [3:0] p15 = (((-2'sd0)?(5'd6):(3'd7))?((-3'sd2)?(5'd18):(5'd8)):((4'd0)?(2'd3):(3'sd0)));
  localparam signed [4:0] p16 = {2{(~(5'sd12))}};
  localparam signed [5:0] p17 = (~&(~|(-3'sd0)));

  assign y0 = (~(|(~|$signed((~^(+(~|(~|(($unsigned((((&(~|(!(~|(~$signed(p9)))))))))))))))))));
  assign y1 = (({1{a0}}|(b1===b2))>((p12<=a3)||{2{b3}}));
  assign y2 = ((2'd1));
  assign y3 = ((a1===b2)&(p8<<<p1));
  assign y4 = $signed(b5);
  assign y5 = (~|p10);
  assign y6 = (({(p8<<b5),(p4<=b3),(-p16)})<{(a0>=a2),((~&p10)),(a4+p1)});
  assign y7 = ((&(p6?p10:p13))?(|(p15?p11:b3)):((|p8)?(-p1):(!p13)));
  assign y8 = (|((4'd2 * a0)?(+a1):(b5?b3:p14)));
  assign y9 = ({1{((b5!==a5))}}^~(&({3{a5}}<<<(p13||a0))));
  assign y10 = (3'd7);
  assign y11 = $unsigned({4{((p6))}});
  assign y12 = ((((b3>>b0)|(a1>=a4))<<((b1|b5)!==(a0<<a1)))&(((a4<<a5)*(a3>>b0))||((6'd2 * a0)!=(a3!=a0))));
  assign y13 = {b4,a1};
  assign y14 = ({1{($unsigned((~b4))^~(b3?a2:b2))}}+((b1?a1:b5)<$unsigned((a3|a5))));
  assign y15 = ((((p13?a2:b3)?(~b3):{b4,a5})<<<{3{(&b1)}})^(~&{(b0?b4:a2),(b4||b3),(p15-p14)}));
  assign y16 = (2'sd0);
  assign y17 = ($signed({(~&(-{3{p5}})),{1{$unsigned({4{a2}})}}}));
endmodule
