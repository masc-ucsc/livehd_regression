module expression_00616(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd1)?(3'sd1):(-5'sd15))?((5'sd3)?(3'sd3):(-4'sd6)):((5'sd14)?(2'd2):(2'd1)));
  localparam [4:0] p1 = ((5'd6)<=(3'd0));
  localparam [5:0] p2 = (~|{(-(((4'd6)?(5'd12):(2'sd1))<<<(2'sd0))),((-3'sd2)?((3'sd3)?(-3'sd2):(2'd3)):((4'd12)?(5'sd14):(-3'sd2)))});
  localparam signed [3:0] p3 = (~^(+(|(~&(~|(&(~&(-(^(^(&(^(&(~|(+(5'd29))))))))))))))));
  localparam signed [4:0] p4 = ({4{((-3'sd0)|(4'd13))}}+(((4'sd6)&&(2'd3))?{3{(5'sd15)}}:((5'd1)<<<(4'sd5))));
  localparam signed [5:0] p5 = {4{{(+((4'sd0)?(4'd8):(2'd2)))}}};
  localparam [3:0] p6 = (2'sd0);
  localparam [4:0] p7 = (+(2'd1));
  localparam [5:0] p8 = ({((3'd2)>=(5'sd14)),{(3'sd3)},((-4'sd4)?(5'sd3):(-3'sd1))}?{((5'd9)?(2'd0):(-3'sd3))}:({(2'd1),(4'sd2),(5'd14)}?{(4'd13)}:{(-5'sd3)}));
  localparam signed [3:0] p9 = {2{((4'sd4)?(-3'sd0):(2'd0))}};
  localparam signed [4:0] p10 = ({2{((5'd31)===(3'sd0))}}===((3'sd2)>>>{(4'd11)}));
  localparam signed [5:0] p11 = (((3'd7)<={3{(3'd2)}})<=(~{(-(4'sd0))}));
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = (4'sd4);
  localparam [5:0] p14 = {{(+(3'sd3)),{3{(2'sd0)}}},(+(^{3{(-4'sd2)}})),(^(&(3'sd2)))};
  localparam signed [3:0] p15 = (5'sd0);
  localparam signed [4:0] p16 = (-2'sd0);
  localparam signed [5:0] p17 = (~&(((5'd16)?(3'd5):(4'd12))?(~((2'd3)?(-3'sd0):(2'd1))):((5'd28)?(5'd9):(2'd1))));

  assign y0 = (&(((a3^a1)===(^a1))^((a1>>>a2)^(b4!=p13))));
  assign y1 = (p4?p4:p15);
  assign y2 = (6'd2 * (p14<<p1));
  assign y3 = (!(p7^~p1));
  assign y4 = (&((~^(5'd1))>>>(3'd3)));
  assign y5 = ($unsigned({({a4}<<(p9|p12))})-{(p5),(a1!==a4),(p6&&p6)});
  assign y6 = ((($unsigned(({a4,b3,a4}!==((6'd2 * b0)||{a5,a1,b3})))==(($unsigned(p3)&{p4})-{(p9&p8),(p13>=p7)}))));
  assign y7 = (~|(+(&p6)));
  assign y8 = (-2'sd0);
  assign y9 = (-4'sd7);
  assign y10 = $unsigned(((4'd1)?$signed($unsigned(b4)):(b3^p6)));
  assign y11 = (4'sd7);
  assign y12 = {{4{p1}},({b5}>>{1{b2}}),(5'd4)};
  assign y13 = ($unsigned($signed((p7>>a1)))==(|(+(+(p2?b2:b5)))));
  assign y14 = $unsigned((-3'sd3));
  assign y15 = {2{{4{(+p14)}}}};
  assign y16 = ((5'd24)!==((4'd10)<<<(b1?a3:a0)));
  assign y17 = {1{(~{({(~^((p14?p1:p10)?{p6}:(p0-p9)))}<(^(-$signed(((p0<<p10))))))})}};
endmodule
