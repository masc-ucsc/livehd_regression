module expression_00671(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^((-5'sd7)||(3'sd1)))%(5'd6));
  localparam [4:0] p1 = (|((~((2'sd0)<(3'sd0)))/(5'd21)));
  localparam [5:0] p2 = (&((((-5'sd14)||(-2'sd0))^~(5'd24))&&(((4'sd4)!==(-2'sd0))==(~^(3'sd1)))));
  localparam signed [3:0] p3 = ((((-2'sd0)>=(5'd5))?((3'd3)+(-3'sd3)):(-5'sd0))<<(((5'd16)?(4'sd0):(5'sd11))>((-3'sd0)^(-4'sd4))));
  localparam signed [4:0] p4 = (^(-2'sd0));
  localparam signed [5:0] p5 = (((4'd0)?(2'd1):(3'd3))?(2'sd0):(4'sd7));
  localparam [3:0] p6 = (3'd5);
  localparam [4:0] p7 = ((~^(3'd3))>>(^(4'd6)));
  localparam [5:0] p8 = {1{((4'sd6)-(5'sd4))}};
  localparam signed [3:0] p9 = (^(-2'sd0));
  localparam signed [4:0] p10 = {(4'd2)};
  localparam signed [5:0] p11 = ((-4'sd3)!==(5'd30));
  localparam [3:0] p12 = (!(((3'd2)===(4'd8))||(4'd2 * (2'd0))));
  localparam [4:0] p13 = (-3'sd1);
  localparam [5:0] p14 = (((!(5'sd8))+(~&(4'sd4)))!==(~{(~|{(-5'sd2),(-3'sd1),(4'd10)})}));
  localparam signed [3:0] p15 = ((2'd3)>(3'd6));
  localparam signed [4:0] p16 = ((5'd1)<<(~^(+(-((4'd14)-(5'sd1))))));
  localparam signed [5:0] p17 = (^(^(~(5'd23))));

  assign y0 = {2{(-2'sd0)}};
  assign y1 = (~^{(~(($unsigned({p8,b4,p15})<(a4!==a4))>>(!((p11)?{1{p14}}:{b4,b3}))))});
  assign y2 = (($unsigned($signed($signed(($unsigned((6'd2 * p6))))))|$signed(((($signed(p3)&&(b5)))))));
  assign y3 = ({2{(3'd4)}}?{3{p8}}:(p2?p1:p9));
  assign y4 = ((p2>p11)^{4{p1}});
  assign y5 = {1{{3{{4{p4}}}}}};
  assign y6 = {2{{{{4{p15}}},{{1{p4}},{2{p12}}}}}};
  assign y7 = ({1{((^{2{p8}})+(5'd7))}}<<(+(2'd3)));
  assign y8 = {4{(|(p3?b1:p10))}};
  assign y9 = ((2'd2)<<$signed(b5));
  assign y10 = ({2{(((b5<b1)>>>(3'd0)))}}!==(((b1<a5)>(b1?a1:b5))&&($unsigned(a4)>{4{a2}})));
  assign y11 = {3{(b5===b3)}};
  assign y12 = {{p0,p0,b0}};
  assign y13 = ((~{3{(p17+p3)}})?((p1>>p8)>>$unsigned((!p7))):{2{$signed((p11^p15))}});
  assign y14 = (-2'sd0);
  assign y15 = $signed((~^($unsigned((5'd14))^((b0<b5)>>>(3'd1)))));
  assign y16 = (((p15?p16:p17)?(~p3):(p12?a3:p3))?(~|((p0?p0:p10)?(p11?p4:p9):(p4==a3))):((p15?p12:p2)<<<(p3&&p17)));
  assign y17 = (b4^~b0);
endmodule
