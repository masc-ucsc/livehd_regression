module expression_00870(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(+((+(-(5'd12)))?((3'd5)?(-4'sd0):(4'sd3)):(5'd2))));
  localparam [4:0] p1 = (~^((((5'd6)!==(-4'sd0))^~((3'd5)?(-4'sd5):(4'd4)))?(((3'sd1)&&(-2'sd0))<=((4'd10)>>(4'd8))):(~^(~(~(+(3'sd1)))))));
  localparam [5:0] p2 = (((-{(3'sd0),(2'd2),(3'd3)})==={3{(5'd29)}})==={4{(&(3'sd1))}});
  localparam signed [3:0] p3 = {{(3'd0)},{(4'd1),(5'sd3),(2'd1)},{(2'd1),(2'sd1),(3'sd1)}};
  localparam signed [4:0] p4 = {((!(-3'sd0))==((4'd6)>=(-2'sd0))),(|({(-3'sd1),(3'd2),(4'd3)}^((-5'sd15)!==(-2'sd0))))};
  localparam signed [5:0] p5 = (4'd11);
  localparam [3:0] p6 = (~(~(2'sd0)));
  localparam [4:0] p7 = ((-5'sd2)?{(5'sd8),((5'sd6)?(4'd9):(4'd14))}:(((-3'sd3)<(5'sd4))+{(2'd1),(3'sd1)}));
  localparam [5:0] p8 = (((3'd5)>=(3'd6))||{(2'd3),(3'd2),(-4'sd0)});
  localparam signed [3:0] p9 = (-5'sd2);
  localparam signed [4:0] p10 = ((+((~^(-3'sd2))!=((5'sd10)<=(5'd20))))<{(^((4'sd6)>>>(4'd10)))});
  localparam signed [5:0] p11 = {{2{(2'd1)}},(~(5'd0)),{1{(4'd7)}}};
  localparam [3:0] p12 = {(!(3'sd3)),(~^(3'd2))};
  localparam [4:0] p13 = ((2'd1)>>>(((-4'sd6)^(3'd2))?((4'sd0)?(3'd6):(4'd14)):(^(5'd17))));
  localparam [5:0] p14 = {(((-5'sd5)<(4'd1))==((2'd3)||(4'sd2))),{((5'sd3)?(2'd2):(4'd6)),((2'sd0)<=(4'sd1)),{(3'sd1),(5'sd13)}}};
  localparam signed [3:0] p15 = {(~^{{(4'd14),(4'sd3),(-5'sd3)},{(2'd2),(2'd0),(4'sd7)}}),(-(!{{(5'd2),(-2'sd1),(5'sd14)},(~^(-2'sd1)),{(5'd11)}}))};
  localparam signed [4:0] p16 = {(3'sd0)};
  localparam signed [5:0] p17 = (5'd8);

  assign y0 = (~^{2{(|(($unsigned((p14<=a2)))))}});
  assign y1 = ({1{((6'd2 * p14)<<(a2+b0))}}&&((b0?a3:b2)?(5'd2 * p8):(b4<=b3)));
  assign y2 = (|((!((p9?p12:p0)?(b1+p4):(~^b5)))?{(-a3),{p2,b5,b3},(+a2)}:((~^p3)?(p4?p16:a5):(b5?p2:p10))));
  assign y3 = $unsigned(({(+(!(b5!=b0)))}?((b5?b0:a2)<<<(~&a5)):(~(6'd2 * (!b1)))));
  assign y4 = ((a1<a3)==(2'd2));
  assign y5 = ({2{$signed($unsigned((b3^~b3)))}}>>>($signed({3{a4}})?$unsigned((a4)):(a0^a1)));
  assign y6 = {1{(&((+(-{4{b3}}))<<<((~p1)>(~b0))))}};
  assign y7 = {(a3&p17),{p13},$signed(p1)};
  assign y8 = (+((b0===b5)<=(b3<=b2)));
  assign y9 = (5'd14);
  assign y10 = ($unsigned((($signed((b3===b5))-{3{p7}}))));
  assign y11 = (-4'sd2);
  assign y12 = $unsigned($unsigned((((-5'sd12)>>(&a1))-{4{a0}})));
  assign y13 = (p8|p11);
  assign y14 = ((p14?p16:p14)?{b0}:(|p9));
  assign y15 = (~^b2);
  assign y16 = (((a1==a2)>=(b0!=p9))+(5'd2 * (p7|b2)));
  assign y17 = (3'd4);
endmodule
