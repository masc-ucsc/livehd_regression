module expression_00234(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~&(-5'sd6))<<<(5'd6));
  localparam [4:0] p1 = (~^({((2'd3)<=(4'd3))}!=((4'd6)?(4'sd7):(-3'sd3))));
  localparam [5:0] p2 = (~(((2'sd1)==(4'sd5))===(|(~^(4'd7)))));
  localparam signed [3:0] p3 = (|(-(&(-(~((2'd1)+(5'd3)))))));
  localparam signed [4:0] p4 = ((5'd19)&(4'sd7));
  localparam signed [5:0] p5 = (~(((2'sd1)<<<(4'sd5))%(5'd15)));
  localparam [3:0] p6 = (^(2'd0));
  localparam [4:0] p7 = (((5'd1)^(-5'sd5))<((4'd15)-(3'd4)));
  localparam [5:0] p8 = ({4{((3'sd1)?(3'sd3):(5'd13))}}>(3'd0));
  localparam signed [3:0] p9 = {1{{1{(2'sd0)}}}};
  localparam signed [4:0] p10 = ((+(-3'sd0))>=((3'sd1)!==(-4'sd7)));
  localparam signed [5:0] p11 = (|((((2'd2)?(-2'sd1):(4'd11))^(~^(5'd23)))||((!(-2'sd1))>=((2'd0)?(5'd27):(-3'sd3)))));
  localparam [3:0] p12 = {2{{1{({4{(2'sd0)}}&&{(2'd3),(5'd21)})}}}};
  localparam [4:0] p13 = (|(^{4{(~|(5'd23))}}));
  localparam [5:0] p14 = {4{{(-4'sd2),(5'd2),(2'sd0)}}};
  localparam signed [3:0] p15 = {((~&(-4'sd2))?((-2'sd0)?(-4'sd7):(5'sd2)):((4'd15)?(4'd8):(-2'sd1))),{{((4'sd6)?(4'd1):(3'd3)),((-4'sd0)?(-5'sd12):(5'd11))}}};
  localparam signed [4:0] p16 = {4{(5'd1)}};
  localparam signed [5:0] p17 = ((((2'd0)?(2'd0):(-5'sd11))?((-4'sd3)<=(-2'sd1)):((2'd0)^~(5'd26)))^(((3'sd2)?(3'd2):(3'sd3))||((3'd7)?(-3'sd1):(4'sd5))));

  assign y0 = (((&(b5))!==(b1||a4))===(4'd4));
  assign y1 = (-((-p13)<(p14<=a4)));
  assign y2 = (-$signed((~$unsigned(((^(~p15)))))));
  assign y3 = (4'd15);
  assign y4 = {$signed({p14,p1,b0}),{p13,p3,p0},$signed($unsigned((2'sd0)))};
  assign y5 = {{$signed(a1),{b5},(b1&&a0)},{(a4-b0),$signed(a0)},((a4^~p5)^~(b5||p16))};
  assign y6 = (((p0&a0)&(a1!==a4))&((p7<<<p8)^(p1<<p2)));
  assign y7 = (p11?p3:p8);
  assign y8 = (3'sd0);
  assign y9 = ({2{(a4|b5)}}>>(4'sd7));
  assign y10 = ({(p16?p16:p7)}?{1{(&(p15>>p4))}}:((!a0)^{p2,p9,p8}));
  assign y11 = (2'd0);
  assign y12 = (!{1{{2{((|{2{b5}})>(~(p12+b2)))}}}});
  assign y13 = {(($signed((b3||b1))>(b1<<<b1))),(~|(6'd2 * (a2-a2))),(((^(b4==b2))===(a5>>a3)))};
  assign y14 = $signed((~{1{b0}}));
  assign y15 = {3{((p2<p14)==(~p3))}};
  assign y16 = ((p6?b4:b3)?((a4&&a5)*(a2?a0:p14)):(4'd0));
  assign y17 = {2{($unsigned((p3>>p7)))}};
endmodule
