module expression_00396(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd1)?(3'd4):(4'd3))>(&(4'sd3)));
  localparam [4:0] p1 = ({(4'sd6),(2'sd1)}|((4'sd3)-(2'd0)));
  localparam [5:0] p2 = ((((-3'sd3)^~(5'd10))-{3{(2'd2)}})?{(3'd1),(-2'sd1),(-3'sd0)}:{{1{((2'd1)?(4'd12):(4'd13))}}});
  localparam signed [3:0] p3 = (((((3'sd2)-(-5'sd9))-((4'd3)<<<(-5'sd3)))+(((2'sd0)>=(3'd7))||((5'd12)<(2'sd1))))&((((4'sd5)-(2'd3))&((3'd1)!=(2'd3)))<=(5'd2 * (2'd1))));
  localparam signed [4:0] p4 = ({(3'd0)}?(2'sd0):(^{((3'sd2)|(5'd29))}));
  localparam signed [5:0] p5 = ((|{3{(5'd25)}})&&(5'd19));
  localparam [3:0] p6 = ((-5'sd1)-(3'd5));
  localparam [4:0] p7 = (-(!{{(-2'sd0),(2'd1)},((2'd2)+(2'd3)),((2'd0)>>(3'sd0))}));
  localparam [5:0] p8 = {4{((-2'sd0)?(-3'sd0):(3'sd3))}};
  localparam signed [3:0] p9 = ((4'd15)===(-4'sd3));
  localparam signed [4:0] p10 = (&{1{((-5'sd0)===(-5'sd13))}});
  localparam signed [5:0] p11 = {2{((3'd7)?(5'd2):(3'sd2))}};
  localparam [3:0] p12 = ((-5'sd4)|(-2'sd0));
  localparam [4:0] p13 = {4{(5'd16)}};
  localparam [5:0] p14 = {((^{4{(2'd2)}})+(|{(~|(4'sd4))}))};
  localparam signed [3:0] p15 = ({((&(!(5'sd15)))>=(&(~|(3'd4))))}+{4{((2'sd0)<=(-3'sd3))}});
  localparam signed [4:0] p16 = {3{(4'sd0)}};
  localparam signed [5:0] p17 = ({((3'd7)<<<(2'd2)),{((5'sd7)&&(2'sd0))}}+({((-4'sd0)|(4'd2))}+((2'd0)>>(2'd3))));

  assign y0 = (((a1<a5)===$unsigned((b0<=b1)))>={4{(b4||b4)}});
  assign y1 = (p3%p10);
  assign y2 = (~&(~|((p4>p12)/p5)));
  assign y3 = $unsigned(($signed((4'd2))&((a2?p10:p14)|((4'sd6)&&(b1&b4)))));
  assign y4 = {2{{2{$unsigned((4'd2 * p14))}}}};
  assign y5 = {((b2?b2:p11)>>>(a3?a3:a2)),((p3<<p0)>>>(b0|b2)),((a1?b2:p16)?(p3==a4):(p4?p3:a3))};
  assign y6 = {(p9<p6),{p3,p1,p3},(p7?p4:p8)};
  assign y7 = (~|p0);
  assign y8 = $signed((((p14<p14)?$unsigned(a0):(p10?p6:b1))?{4{p4}}:(!(2'd0))));
  assign y9 = ((b3?b3:a4)!==(a4>=b4));
  assign y10 = (&(|(~&a4)));
  assign y11 = ({(~|a0),(a1>>a3),(~&a3)}^~(~^((~&{b4})||{2{p9}})));
  assign y12 = ((b1?b2:a3)%a0);
  assign y13 = (4'd5);
  assign y14 = {4{({3{p1}}>>>(~&a5))}};
  assign y15 = ((|(((-5'sd15)&&{b3,p15})&&{b3,p14,p10}))>{(+(~b5)),(-5'sd4),{a5,p11,p4}});
  assign y16 = ((~(p6|a1))^~{2{(~|a5)}});
  assign y17 = $signed($signed(((5'd16)?(~(2'sd0)):{2{{b2,a2}}})));
endmodule
