module expression_00462(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(~{(!((2'd2)<<(4'd13))),({3{(-5'sd1)}}<<<{1{(3'd0)}}),{1{(-(!(2'd2)))}}})}};
  localparam [4:0] p1 = (^(&(~(~&(~&(+(!(|(+(^(~^(^(&(4'd0))))))))))))));
  localparam [5:0] p2 = ((((5'sd7)>>>(4'sd0))?(!(2'sd1)):((2'd1)?(2'd1):(5'd13)))==(~&((-(&(-2'sd0)))!==(|((2'sd0)===(2'd1))))));
  localparam signed [3:0] p3 = (((~|(3'd7))?((2'sd0)?(2'd0):(3'd0)):(+(3'sd0)))<({(4'd12)}?((4'sd4)?(-5'sd15):(-2'sd1)):(5'd2 * (3'd2))));
  localparam signed [4:0] p4 = {1{(3'd5)}};
  localparam signed [5:0] p5 = ({1{(-2'sd0)}}^(6'd2 * (4'd4)));
  localparam [3:0] p6 = ((|(-3'sd0))||(&(3'sd1)));
  localparam [4:0] p7 = (((^((2'd2)|(3'd3)))/(-3'sd3))|(&(((2'sd0)^~(2'd2))<<<(-(-(2'd3))))));
  localparam [5:0] p8 = {1{({((4'd14)?(-5'sd14):(4'd1)),{1{(3'd1)}},(-(5'd14))}>{2{((2'd1)^~(4'd3))}})}};
  localparam signed [3:0] p9 = ((((2'd1)<=(4'd4))===((3'sd1)^~(3'sd0)))!==(~|{4{(-2'sd1)}}));
  localparam signed [4:0] p10 = (&((~((-2'sd1)^~(3'd6)))?(~&(4'd2)):(4'sd7)));
  localparam signed [5:0] p11 = (~|(-(-(~|(~|(&(~&(~(~^(!(~|(&(3'd2)))))))))))));
  localparam [3:0] p12 = (({(3'd3),(-2'sd0),(2'sd1)}>>>(~&{(-2'sd1),(5'd25),(2'd0)}))+(((3'sd2)?(3'sd3):(3'sd1))>>((5'd14)?(3'd5):(3'sd2))));
  localparam [4:0] p13 = (((-2'sd0)%(3'sd1))?((2'd3)>>(-3'sd2)):(~&(-3'sd3)));
  localparam [5:0] p14 = (((-4'sd5)?(3'sd3):(5'd0))+(!(4'sd5)));
  localparam signed [3:0] p15 = {1{(&(|(-5'sd7)))}};
  localparam signed [4:0] p16 = (((~(4'd14))?(!(4'd7)):((3'sd0)&&(-4'sd3)))?({4{(-5'sd4)}}^((-5'sd0)?(3'd3):(-2'sd1))):(~(|{3{(3'sd1)}})));
  localparam signed [5:0] p17 = {4{(3'sd1)}};

  assign y0 = {1{(&b1)}};
  assign y1 = ((~&(~^(a1?p1:b1)))?(~((-b4)?(p8==b4):(a5===a3))):((a4>>p3)!=(b0?b5:b1)));
  assign y2 = {3{{2{(-{2{a5}})}}}};
  assign y3 = (~(-((~^{2{p1}})||(5'd2 * {1{a1}}))));
  assign y4 = (p9>>>p14);
  assign y5 = (($unsigned(a2)<=(a1+a4))&&({p13,b0,b4}||(+a5)));
  assign y6 = ((~(5'd2 * (b1===b2)))<(4'd7));
  assign y7 = ((~|(!(((!p12)+(p12==b0))<<<(!(a0<<p11)))))!=(&((a0===b1)?(p9^~a2):(2'd3))));
  assign y8 = (5'sd1);
  assign y9 = ((&((a5+b5)?(b1?b2:b3):{b1,a5,b4}))!==(~^(({b2}<<(b0?b0:b1))<<({b2,a0}===(&a5)))));
  assign y10 = (-3'sd2);
  assign y11 = (({1{p17}}=={4{a0}}));
  assign y12 = (((a4?p17:p10)?(b2%a0):(a4>>a4))|((a1?b5:p12)*(p3%b1)));
  assign y13 = {4{(b0<=p3)}};
  assign y14 = (((^(^(b3===b3)))>=((&b4)*(^a5)))^~((~|(~(5'd2 * b1)))==(-3'sd2)));
  assign y15 = $signed({1{(+({4{p13}}>(-{3{p11}})))}});
  assign y16 = (((~&(~&(b4>=a1)))^~((b0||p11)^(~&b2)))^~(+{2{{2{p10}}}}));
  assign y17 = ((~$signed((2'sd0)))?(4'd2 * (!b2)):(+(-5'sd14)));
endmodule
