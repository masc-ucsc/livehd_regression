module expression_00199(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|{3{(+(4'd5))}});
  localparam [4:0] p1 = {{(2'd0),(5'd15)},((3'd4)?(4'sd0):(-3'sd1)),(~(&(3'd7)))};
  localparam [5:0] p2 = (-(3'd1));
  localparam signed [3:0] p3 = (+(-({3{(~^(-5'sd5))}}<(((3'd0)<(5'd7))?((4'd15)<<(4'sd4)):{4{(4'd6)}}))));
  localparam signed [4:0] p4 = {(3'd7),(~^(~^(~&(-3'sd0)))),{(-2'sd1),(-(-4'sd1))}};
  localparam signed [5:0] p5 = (((-4'sd6)?(5'd11):(4'sd4))?(-((-3'sd3)?(-4'sd0):(2'd2))):((3'sd2)?(2'sd0):(4'sd6)));
  localparam [3:0] p6 = (+(|((3'd5)?(5'sd3):(4'd1))));
  localparam [4:0] p7 = ((5'd16)>=(~|(5'd0)));
  localparam [5:0] p8 = (-3'sd0);
  localparam signed [3:0] p9 = ((-2'sd0)^(4'd3));
  localparam signed [4:0] p10 = (-(~^(&(&(|(|(+(-(2'd2)))))))));
  localparam signed [5:0] p11 = (5'd19);
  localparam [3:0] p12 = (~&(^(|(|(|((4'sd3)<<<(3'sd1)))))));
  localparam [4:0] p13 = (-4'sd2);
  localparam [5:0] p14 = (+{4{((-5'sd7)^(5'd23))}});
  localparam signed [3:0] p15 = (&(2'd0));
  localparam signed [4:0] p16 = ((3'd7)?(5'd12):(4'd0));
  localparam signed [5:0] p17 = {1{(5'sd14)}};

  assign y0 = (~&{4{(a3?a3:a5)}});
  assign y1 = (5'd27);
  assign y2 = ({{(p2?a1:b5),(b0?p1:a0)}}?((a3?b2:p0)?{a5,b3,p13}:{p8,p2,a4}):(-2'sd1));
  assign y3 = (((p3?p16:p5)?{3{p0}}:{p8,p7})?({1{{4{a1}}}}+{p3,p12,a3}):{3{{4{p17}}}});
  assign y4 = ($unsigned(((a4-b4)&&{4{a5}}))^{1{((-(a3+p1)))}});
  assign y5 = $unsigned((($unsigned(b2)?(p1>b4):(p15^a1))>(4'd11)));
  assign y6 = (^(((p8>=b2)&&(p1>>>p1))>=({b5,p11}&(a1||a4))));
  assign y7 = $signed({2{(($unsigned((p15<<<a5))==({4{p3}}<$signed(p13))))}});
  assign y8 = (((p7+b0)&&{1{(b2|a5)}})<={3{(p13<a0)}});
  assign y9 = ({(4'd2 * (^(2'd0)))}?{2{{4{p16}}}}:($unsigned((b5!==b2))<<{3{p14}}));
  assign y10 = (((a3?a0:a3)<<{b2})<((b2+b1)==(b4<a5)));
  assign y11 = {(-(~{(&{a5,b1}),{p4,b1,b5},(|{a1,a1,a2})}))};
  assign y12 = (~&(a0^~b1));
  assign y13 = {{(p15&&a3),(~&p15),{p8,p14,p15}},{(~{((5'd2 * p13)<={p14,p8})})},((a0||b2)!==(b3<b4))};
  assign y14 = ({1{(-a3)}}>(b3?p5:b1));
  assign y15 = ((5'd22)<(((5'sd10))<=(-2'sd1)));
  assign y16 = ((a5&b4)%a4);
  assign y17 = (~&{1{(!a5)}});
endmodule
