module expression_00937(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((5'd28)>>(4'd12))^~(4'd7)),{3{(3'd0)}}};
  localparam [4:0] p1 = ((~(4'sd0))?((-3'sd1)==(4'd4)):(~^(4'sd5)));
  localparam [5:0] p2 = (~^(((3'd0)<<(-2'sd0))=={1{((-2'sd1)!==(-4'sd3))}}));
  localparam signed [3:0] p3 = (((((-3'sd3)-(3'd3))^((3'd5)>(2'd1)))&(((4'd13)^~(-2'sd1))<<((-4'sd2)<(4'd15))))>>((((5'sd14)!=(4'd7))<=((-2'sd0)<(4'sd0)))<=(((-2'sd1)^(4'sd7))>((-3'sd3)<<(2'd1)))));
  localparam signed [4:0] p4 = ((-2'sd1)?(5'sd3):(3'sd1));
  localparam signed [5:0] p5 = ({2{((5'd14)+(4'd2))}}-({2{(2'd1)}}?((3'd7)&&(-5'sd14)):((3'd1)^(2'sd0))));
  localparam [3:0] p6 = (((3'sd3)?(-2'sd0):(-4'sd5))-(-3'sd2));
  localparam [4:0] p7 = {1{(-((5'd4)?(3'sd3):(4'sd2)))}};
  localparam [5:0] p8 = (^((~{(3'sd0),(2'sd1),(-4'sd2)})!=(|((4'sd7)-(!(3'd3))))));
  localparam signed [3:0] p9 = {4{((-4'sd0)||(-2'sd0))}};
  localparam signed [4:0] p10 = ((^(5'd26))>(4'd2 * (2'd2)));
  localparam signed [5:0] p11 = (2'sd1);
  localparam [3:0] p12 = (((4'd12)?(2'd0):(-3'sd0))?((2'sd0)+(3'd6)):((5'sd9)==(2'd0)));
  localparam [4:0] p13 = ({(2'sd1),(5'd5),(-3'sd1)}?{(4'd2),(3'd0),(3'sd3)}:(((4'd2)?(3'sd3):(-5'sd2))<((-5'sd10)&(5'd30))));
  localparam [5:0] p14 = (((4'd5)!=(2'sd1))||(^(5'd30)));
  localparam signed [3:0] p15 = (-(~((^(-((~^(2'd3))<((4'sd6)|(4'd7)))))^~(((3'd7)-(4'sd3))||((2'sd0)!==(2'd1))))));
  localparam signed [4:0] p16 = (!(&(~&(((3'sd0)^(3'd7))<(~^(2'sd1))))));
  localparam signed [5:0] p17 = (-3'sd1);

  assign y0 = (((3'sd0)^~(|(4'sd2)))?(((a0<=p5)&&(!(2'd3)))):({a0,p8,a0}+$unsigned({p7})));
  assign y1 = (&((3'd4)!==((a1?a0:a0)>(a5<<a2))));
  assign y2 = ((|(+($signed((+((p5<=p8)&&(b2||b1))))>>$signed((((b2)==(|a2))!==$unsigned((a5|a3))))))));
  assign y3 = {((3'd0)!=(-2'sd1))};
  assign y4 = {3{(+((3'd1)==(p1?a0:p16)))}};
  assign y5 = {3{((!b5)?(b2?p16:b2):(b5===a1))}};
  assign y6 = ({(b4+a1),(a2<b4),(|(~^b4))}^~(((4'd9)>(b2<<<b3))+{b2,b2,a3}));
  assign y7 = $unsigned(p6);
  assign y8 = ((|(5'd1))|($unsigned((3'd7))));
  assign y9 = ($signed(({1{(b0==b2)}}))||{4{{1{a0}}}});
  assign y10 = {3{p9}};
  assign y11 = (!(((b2!==a2)>=(~^p1))?((6'd2 * b2)>=(p9?p3:p1)):({3{p11}}&&(p1-p7))));
  assign y12 = (a1>p5);
  assign y13 = (4'd2 * {2{p13}});
  assign y14 = (4'd2 * (p8==p2));
  assign y15 = {{(a0?b0:p1),(~&{b0,b0,a0})},(2'd0)};
  assign y16 = (+(^{2{a2}}));
  assign y17 = (^((p17>p4)||(2'd2)));
endmodule
