module expression_00384(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd2)?(3'sd2):(3'sd0))?((-5'sd14)<(-4'sd3)):((3'd6)!==(-2'sd0)));
  localparam [4:0] p1 = (-5'sd2);
  localparam [5:0] p2 = (~|({2{(4'sd6)}}>>>(6'd2 * (2'd3))));
  localparam signed [3:0] p3 = (-(2'sd1));
  localparam signed [4:0] p4 = (|((~|((2'd0)?(4'd9):(3'sd3)))?(((-3'sd0)<=(5'd30))!==((5'd28)?(3'sd1):(-4'sd7))):(((-3'sd2)>>>(4'd8))+(!(-2'sd0)))));
  localparam signed [5:0] p5 = {2{(~&(^(~(~&(~^{4{(4'sd7)}})))))}};
  localparam [3:0] p6 = {2{{4{(~(-3'sd0))}}}};
  localparam [4:0] p7 = ((-3'sd1)?(-4'sd0):(2'd3));
  localparam [5:0] p8 = {2{{(2'd1),(4'd13),(-5'sd7)}}};
  localparam signed [3:0] p9 = {2{(5'd12)}};
  localparam signed [4:0] p10 = {2{((5'd0)<<<(2'd1))}};
  localparam signed [5:0] p11 = (~(((-3'sd2)&(4'd9))|(4'd2 * (4'd5))));
  localparam [3:0] p12 = (((4'sd4)>=(-2'sd1))>=(~&((-3'sd0)>>(3'sd1))));
  localparam [4:0] p13 = ({(5'd1),(3'sd1)}&((3'd6)==(3'sd3)));
  localparam [5:0] p14 = (~|(~((((2'd0)*(-5'sd0))<<(4'd2 * (5'd28)))===(((5'sd0)<=(2'd2))*(^(5'sd4))))));
  localparam signed [3:0] p15 = {4{(-5'sd4)}};
  localparam signed [4:0] p16 = ((~&((4'sd3)-(5'd5)))^~(~&(-((3'sd3)?(3'd7):(-5'sd7)))));
  localparam signed [5:0] p17 = (~|(((~&((-3'sd0)!=(5'd4)))==(~(~|(5'sd7))))<(~(~&(((2'd0)*(3'd6))|((4'sd7)&(-5'sd14)))))));

  assign y0 = {3{((p5&p1)-(~&a0))}};
  assign y1 = (a3?a5:a3);
  assign y2 = $unsigned(({a1,p14}?$unsigned({p16,p12}):{p16,b4,p11}));
  assign y3 = (a5-a0);
  assign y4 = (((-b0)?(~|b1):(|b4))?(~(p4?a1:b1)):((-p15)?(~&a1):(&a5)));
  assign y5 = $signed(((2'd2)|((p4^a2)|(5'd11))));
  assign y6 = ((b0?a5:b1)?(p6?p9:b3):(b5?p15:a2));
  assign y7 = ((|((p11^p10)<(p11/p4)))+((a5?b1:a0)===(|(a5>>>b3))));
  assign y8 = (~((!{(!((2'd1)))})-(|$unsigned({2{(3'sd3)}}))));
  assign y9 = (~{3{(3'd3)}});
  assign y10 = {3{a2}};
  assign y11 = {(b2==b3),{b5,p13},{p5,p16}};
  assign y12 = ((^(~(5'd30)))>>>((~{(-p2),(p14>=p7)})<<<{3{{b1,p2}}}));
  assign y13 = ((!$unsigned((4'sd2)))<((~|{p17,p15})&&$unsigned({p13,p7,p6})));
  assign y14 = (~^(-3'sd1));
  assign y15 = ({3{a4}}>=(p13>a4));
  assign y16 = (((a4!=a5)>>>(5'd2 * p13))?((b3>=a2)<<(b5>=p4)):((-2'sd0)&(p5<p0)));
  assign y17 = ((~({p5})));
endmodule
