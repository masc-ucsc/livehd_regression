module expression_00530(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((5'd4)+(-4'sd1))?{(4'd11),(-5'sd14),(2'sd1)}:(~(2'd2))),{1{{{1{{(3'sd1),(4'd9),(-2'sd1)}}}}}}};
  localparam [4:0] p1 = {4{((4'd5)<=(-3'sd3))}};
  localparam [5:0] p2 = (~((3'd2)?(2'd2):(4'sd2)));
  localparam signed [3:0] p3 = (4'd2 * (3'd7));
  localparam signed [4:0] p4 = (({1{(4'sd2)}}?((4'd13)&&(3'sd1)):{4{(-3'sd2)}})||(((-4'sd6)===(-3'sd0))==={(5'sd2),(-2'sd1)}));
  localparam signed [5:0] p5 = ((~(2'd2))<<((4'd12)!==(5'sd10)));
  localparam [3:0] p6 = {{(-3'sd2),(5'd22),(3'sd1)},(^{(4'd7)}),(-(+(5'sd15)))};
  localparam [4:0] p7 = ((+((-4'sd5)&&(2'd1)))?((4'd15)!=(5'd10)):((-4'sd0)%(5'sd5)));
  localparam [5:0] p8 = {4{(5'sd10)}};
  localparam signed [3:0] p9 = (-4'sd3);
  localparam signed [4:0] p10 = (~|(4'd8));
  localparam signed [5:0] p11 = (((5'd2)?(3'd5):(2'sd1))/(3'd0));
  localparam [3:0] p12 = ({((5'd31)?(3'd0):(-3'sd3))}?{((-5'sd12)?(-3'sd3):(2'sd1))}:{(-5'sd14),(-2'sd1)});
  localparam [4:0] p13 = (5'd16);
  localparam [5:0] p14 = ((2'd3)&&({(3'd0),(4'd2),(5'd18)}||((5'd17)^(-4'sd2))));
  localparam signed [3:0] p15 = (~^(!(~&(!{(3'sd0),(4'd10)}))));
  localparam signed [4:0] p16 = (3'd5);
  localparam signed [5:0] p17 = (((3'd6)^(3'd3))<{3{(5'd28)}});

  assign y0 = (|(~^(|((~&(~((!(~&p3))<(~|(p3+a4)))))>>>(-4'sd1)))));
  assign y1 = ((a1-p15)?(-2'sd1):{2{p7}});
  assign y2 = {1{(((b1^~b5)===(-4'sd4))|(&{p14,a3,p4}))}};
  assign y3 = {(|({b5,a5}^(|(!a1))))};
  assign y4 = {2{(a1!==b2)}};
  assign y5 = (4'sd0);
  assign y6 = (((a2>a5)<={3{b3}})!==(&(a1!=a3)));
  assign y7 = {4{((b5?b0:p3)<<<(p6>p8))}};
  assign y8 = $signed($signed({3{$unsigned(p6)}}));
  assign y9 = ($unsigned(p0)-(~^a2));
  assign y10 = (6'd2 * {3{p0}});
  assign y11 = ((b2&&a3)===(a4!=a5));
  assign y12 = (~({(p10?b5:p13)}?(+{1{(p12?b1:b1)}}):(!{3{p9}})));
  assign y13 = (^(^(~^(|(+(((p1)?(+p0):(-p1))?(~|((b5<<<p6)&&(a4?p5:a1))):(~&(~((a3?p2:p14))))))))));
  assign y14 = {($unsigned((-3'sd1))!==$unsigned($signed(a2))),(((b2===b2)>=(-5'sd9)))};
  assign y15 = (((p11/p7)>(^p9))|((~p16)/p13));
  assign y16 = {1{(^{2{({(~(~(^(~^(!(|p2))))))})}})}};
  assign y17 = ((~|$unsigned($signed((|(-2'sd1))))));
endmodule
