module expression_00033(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd7);
  localparam [4:0] p1 = ((((5'd19)-(-2'sd1))&(~&((-3'sd1)>>(-2'sd1))))!==(5'd2 * ((4'd13)<(2'd1))));
  localparam [5:0] p2 = {((-3'sd3)?(4'd9):(4'd10))};
  localparam signed [3:0] p3 = ({(-2'sd0),(3'sd0),(3'd2)}!==((2'd1)+(4'sd0)));
  localparam signed [4:0] p4 = ((4'd15)!==(&{4{{2{(-3'sd3)}}}}));
  localparam signed [5:0] p5 = {(((5'sd0)<<(4'd0))!=((4'd8)!==(2'd3))),(3'd1),(&((+(2'sd1))<{(-3'sd0),(4'd13),(-2'sd1)}))};
  localparam [3:0] p6 = ((((3'sd0)?(3'sd3):(5'd7))?(4'd2 * (5'd6)):(-5'sd6))?(~&((5'd18)?(2'sd0):(2'd1))):((5'd6)||{4{(3'd7)}}));
  localparam [4:0] p7 = {((3'sd3)<(4'sd5))};
  localparam [5:0] p8 = ((~^(-4'sd6))<=(-(-3'sd1)));
  localparam signed [3:0] p9 = {2{{4{(2'sd1)}}}};
  localparam signed [4:0] p10 = (4'sd2);
  localparam signed [5:0] p11 = (~&{(4'd10)});
  localparam [3:0] p12 = {1{{{{(4'd4),(2'sd0)},(!(3'sd0)),((5'd18)<(4'd6))},{(~^(-5'sd13)),{(2'd0),(5'sd8)}},(5'd2 * {1{(|(2'd1))}})}}};
  localparam [4:0] p13 = {(4'd5),(2'd3),(2'd0)};
  localparam [5:0] p14 = (-{{(5'd15),(3'd0),(2'd1)},((4'd12)?(5'd24):(-2'sd0)),((5'd26)?(-5'sd9):(4'd8))});
  localparam signed [3:0] p15 = (5'd6);
  localparam signed [4:0] p16 = {2{(4'sd6)}};
  localparam signed [5:0] p17 = (~|(-(4'd3)));

  assign y0 = (3'd2);
  assign y1 = (+{1{$signed({2{(|(-4'sd0))}})}});
  assign y2 = (4'd3);
  assign y3 = ($unsigned((!(4'd8)))<=(~|(-(b2?p7:b4))));
  assign y4 = $unsigned({1{((~|(p10&&b0))^~((p17|a0)))}});
  assign y5 = (!p8);
  assign y6 = ((p0?p7:p12)?(a4?a5:p0):(p9?a2:p13));
  assign y7 = (~|((3'd2)<(5'd27)));
  assign y8 = ({2{(p15-p3)}}<=(2'd0));
  assign y9 = ((p2-p1)*(p2-p0));
  assign y10 = (+(-(a1*a5)));
  assign y11 = (3'sd0);
  assign y12 = ((b0+a4)^{a4,b2});
  assign y13 = ((|$signed(a5))<(b4?b5:a1));
  assign y14 = (((~&(($signed(p7)^~$unsigned(p14)))))||{3{(b3)}});
  assign y15 = (~^((a5?a4:b0)?((a3?b4:a2)<<{3{b3}}):((|(b1)))));
  assign y16 = (b2?b3:a5);
  assign y17 = {(|$unsigned((4'sd0))),(~|(4'd2 * (a2>=b2)))};
endmodule
