module expression_00925(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-3'sd2)>(-4'sd5))!==((5'd6)>>(5'd2)));
  localparam [4:0] p1 = (~|{4{((-3'sd0)&&(2'd3))}});
  localparam [5:0] p2 = (+((-3'sd0)^~(3'd3)));
  localparam signed [3:0] p3 = (|(~^{(|{(5'd15)}),{(-(2'd0))}}));
  localparam signed [4:0] p4 = {1{({2{{(5'd3)}}}-{({(-4'sd4)}||((2'sd1)>(-3'sd0)))})}};
  localparam signed [5:0] p5 = (|(~|({3{(5'sd5)}}>>>((4'sd7)<(-4'sd5)))));
  localparam [3:0] p6 = ((((5'd12)?(-3'sd2):(5'd15))==((3'd0)&&(5'd17)))?(~&(!{3{(-2'sd1)}})):(!((-2'sd1)?(4'sd4):(-5'sd4))));
  localparam [4:0] p7 = (5'd28);
  localparam [5:0] p8 = (3'sd0);
  localparam signed [3:0] p9 = {4{((-4'sd6)!==(5'sd10))}};
  localparam signed [4:0] p10 = ((6'd2 * (5'd30))?{2{(5'd24)}}:((3'd2)&&(-2'sd0)));
  localparam signed [5:0] p11 = (((4'd6)?(-4'sd0):(-5'sd14))>=(~^{3{(4'd3)}}));
  localparam [3:0] p12 = (((-3'sd1)&(-2'sd0))>=((3'sd0)<=(-2'sd0)));
  localparam [4:0] p13 = (4'sd4);
  localparam [5:0] p14 = (({(3'd0),(4'd2),(4'sd2)}<<{(5'd8),(2'd2)})^(~^({(2'd1),(2'sd1),(2'd1)}!=((-5'sd12)==(2'd3)))));
  localparam signed [3:0] p15 = {3{{4{(5'd18)}}}};
  localparam signed [4:0] p16 = ({3{(-2'sd0)}}&((6'd2 * (3'd7))<=((3'd1)-(2'sd1))));
  localparam signed [5:0] p17 = (&{{{(-(~^{(2'd0)})),(~|{(|(3'sd0))})}}});

  assign y0 = ((((b1<<p0)>>>(p16>>p3))!=$unsigned((!(|a5))))>=(!(&$unsigned($unsigned($signed((p10<p17)))))));
  assign y1 = (((~|((b5!=a0)^~(p9>p3)))!=(-(-(p11<a1))))<<(((b3>>p15)^~(p9-p9))<((a0!==b5)<<<(p5<<<p10))));
  assign y2 = {4{{4{p11}}}};
  assign y3 = (&(5'd2 * (p6&&p6)));
  assign y4 = {1{(p12<p3)}};
  assign y5 = (2'd1);
  assign y6 = {1{{4{(4'sd3)}}}};
  assign y7 = (((~|p2)?(2'sd0):(|a5))?((a2?a3:b5)===(^(~|a4))):(4'd3));
  assign y8 = $signed(((!{1{(+(~^b0))}})));
  assign y9 = (-({b2,b1}>>(|(~^b0))));
  assign y10 = {(^(~(({b1,b1,b5}>>$signed(p8))?{$signed({1{p8}})}:($unsigned(b2)>={2{p15}}))))};
  assign y11 = $unsigned((((3'd3)<=((b0?p11:p11)>>(5'd6)))));
  assign y12 = (~(|{1{{3{{3{p0}}}}}}));
  assign y13 = (-(~|$signed($signed(p1))));
  assign y14 = {(~&((((a4<<p1)&$signed(p12))?(-(b0===a0)):((6'd2 * p7)<<{p8,b3}))))};
  assign y15 = $unsigned(({3{(a1===b1)}}>={4{(b4<<a3)}}));
  assign y16 = {a4,b0,b3};
  assign y17 = {4{(3'd3)}};
endmodule
