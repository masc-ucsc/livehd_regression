module expression_00978(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{{3{{(-2'sd1),(5'sd13)}}}}};
  localparam [4:0] p1 = (!((6'd2 * {2{(5'd0)}})<={2{(~(5'd7))}}));
  localparam [5:0] p2 = ((5'd6)?(&(-2'sd1)):(5'sd13));
  localparam signed [3:0] p3 = (-4'sd2);
  localparam signed [4:0] p4 = {{{{(-3'sd0),(5'sd10),(5'sd2)},((5'd12)^~(4'd8))},(((4'sd0)>>>(2'd1))-{(3'd6)}),{(-4'sd0),(4'd10),(5'sd9)}}};
  localparam signed [5:0] p5 = {3{{(-5'sd7),(3'd7)}}};
  localparam [3:0] p6 = (-4'sd4);
  localparam [4:0] p7 = ({(5'd0),(3'd1),(-2'sd0)}^((2'd1)<<(3'd7)));
  localparam [5:0] p8 = ((3'd4)>>>(2'd3));
  localparam signed [3:0] p9 = ((+((-5'sd11)&&(4'd15)))&&(((5'd12)<<(5'd24))==((2'sd0)%(3'd7))));
  localparam signed [4:0] p10 = (((3'd7)?(4'd8):(-2'sd0))?(&((4'sd6)!=(5'sd8))):{((5'sd1)||(5'd2)),(5'd24)});
  localparam signed [5:0] p11 = (6'd2 * (~|(4'd2 * (3'd3))));
  localparam [3:0] p12 = (~&(~^((&(~&(~(+(&(-2'sd1))))))^~(((4'd1)*(3'sd1))+((3'sd2)<<<(5'd20))))));
  localparam [4:0] p13 = {(3'd7),(2'sd0)};
  localparam [5:0] p14 = ((5'd8)^(~(5'd15)));
  localparam signed [3:0] p15 = {4{(^(~&(3'd4)))}};
  localparam signed [4:0] p16 = (!((|(~^(5'sd11)))||{3{(-2'sd1)}}));
  localparam signed [5:0] p17 = {2{(-3'sd2)}};

  assign y0 = (~^{{((b0<<<p3)?(~&a3):{a3,p8,a4}),((p16!=p10)?{p3,p12,p1}:(~p13))}});
  assign y1 = ({$signed(b4),$signed(a0),(b3|a0)}<<($signed(a0)?(a0&&a0):(p17?b1:a0)));
  assign y2 = ((a1>>a0)/a2);
  assign y3 = $unsigned((p7<p16));
  assign y4 = (b1<<<b4);
  assign y5 = (~&{(-(-{4{p6}}))});
  assign y6 = ((&((a2<<<p12)?(~^p0):(b2<<<p17)))|(!((b2^b2)>>(|p4))));
  assign y7 = (((a0>=a1)<<<{a5,b1,a3})^~({4{b3}}&{(a1==p2)}));
  assign y8 = (-4'sd7);
  assign y9 = (p17);
  assign y10 = (5'd25);
  assign y11 = (-3'sd2);
  assign y12 = ((b0^a4)?(~(b0<a4)):{a4,p8,b3});
  assign y13 = ((((p12&&a1)>>(a0))^~((b3-b0)<=(b2)))<<$unsigned((((a3+b3)!==$signed(b1))&((b4/a2)^(b4/b3)))));
  assign y14 = {3{(5'sd4)}};
  assign y15 = (-(-4'sd5));
  assign y16 = {4{p1}};
  assign y17 = (~|(+((-((~b0)?$unsigned(b1):(b1))))));
endmodule
