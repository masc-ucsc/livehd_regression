module expression_00330(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd1);
  localparam [4:0] p1 = {1{{(2'd2)}}};
  localparam [5:0] p2 = (5'sd11);
  localparam signed [3:0] p3 = ((4'd1)|((&(4'd3))>={3{(2'd2)}}));
  localparam signed [4:0] p4 = (~|((~|((2'd1)<=(5'd24)))<(~^((5'd4)<<(3'd1)))));
  localparam signed [5:0] p5 = ((~(2'sd1))?(((2'd3)&&(4'sd2))<<((4'd1)?(-3'sd0):(5'd28))):(((2'd1)?(4'd7):(-5'sd10))<<<(5'd2 * (5'd7))));
  localparam [3:0] p6 = {1{(3'd6)}};
  localparam [4:0] p7 = ((!{2{((2'd1)==(-3'sd2))}})?((+(-2'sd1))?((-4'sd3)?(5'd22):(4'sd7)):(&(-3'sd1))):((~(5'sd9))?{3{(5'sd6)}}:(~(5'sd11))));
  localparam [5:0] p8 = ((2'd0)?(2'd0):(-3'sd1));
  localparam signed [3:0] p9 = {2{(^({3{(3'sd2)}}==={(2'sd1),(-4'sd3)}))}};
  localparam signed [4:0] p10 = (~|((2'd2)<(5'sd3)));
  localparam signed [5:0] p11 = {1{{4{((5'd22)?(2'd1):(-3'sd2))}}}};
  localparam [3:0] p12 = ((5'd3)>=(&(((2'sd1)/(5'sd11))/(4'd10))));
  localparam [4:0] p13 = {(-5'sd8),(4'sd2),{1{(+((5'd24)>>(-4'sd0)))}}};
  localparam [5:0] p14 = (4'd1);
  localparam signed [3:0] p15 = ((~{3{(4'd7)}})&(!((~(2'd2))^~(3'd1))));
  localparam signed [4:0] p16 = (~(((3'd7)>>((2'd2)>>(-2'sd1)))>>((2'd1)?(2'd2):(2'd1))));
  localparam signed [5:0] p17 = (~&{1{{1{(4'd4)}}}});

  assign y0 = ((5'd17)|(((a0||b1)-(a4<=a2))^~({p12,b2,b2}>(b5?b0:a0))));
  assign y1 = (((a0?p12:p5)?{3{p13}}:(p2?p10:p1))?((p0-p17)>>>$signed((~^p5))):(~((~^p0)||{4{p8}})));
  assign y2 = $signed($unsigned(({1{a4}}===(b3))));
  assign y3 = (-3'sd0);
  assign y4 = (5'd6);
  assign y5 = (((~p17)-(p4>>>p13))||((a0==p4)<<(a3==p12)));
  assign y6 = ((~^(5'd14))?(5'd12):((-4'sd2)+(&b0)));
  assign y7 = (^(((p8<=p8)>(b4))));
  assign y8 = {{(a0^a4),(p15-p3),(p6>>p16)}};
  assign y9 = ((~&({4{b4}}>=(-4'sd6)))<((a4?b2:a3)!==(a3?b1:b5)));
  assign y10 = (^{(a4>=b4),(p10>>p10),(+p4)});
  assign y11 = {($unsigned((p2|b2))<<({p14,a3}|$unsigned(p17))),(((b0!==b4)&(-4'sd6))||(5'sd6))};
  assign y12 = ($unsigned((p1|p7))&&{b0,b1,b5});
  assign y13 = {3{b1}};
  assign y14 = (&(~^({3{{2{a3}}}}^~(&(-(~|(~&{2{b0}})))))));
  assign y15 = $unsigned((((p6)?(p5?p15:p5):(p14-p13))<<(6'd2 * (p12-p6))));
  assign y16 = ({4{a0}}-(p8<=p0));
  assign y17 = $unsigned(((^$signed(($signed((b4!==a3))+(4'd2 * $unsigned(p14)))))+(+(((p11!=a2)==(b1<<<a5))>(-(~^$unsigned(a2)))))));
endmodule
