module expression_00516(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({{(-2'sd0),(5'sd6)},{(3'sd2),(4'd14),(3'd0)},{(3'sd2),(-4'sd5)}}==(((4'sd1)<<(2'd2))==={(4'sd0),(4'sd5),(-2'sd0)}));
  localparam [4:0] p1 = (((5'sd2)-(5'sd0))===(+(^(5'd15))));
  localparam [5:0] p2 = (~&(2'd3));
  localparam signed [3:0] p3 = (({(-5'sd7),(2'sd1)}<{(4'd2)})?(((2'd0)<<<(2'd3))?((5'd1)?(4'd11):(5'd2)):((2'd3)<<<(-2'sd0))):{{4{(3'd3)}}});
  localparam signed [4:0] p4 = (&(((-5'sd12)*(3'd1))?((2'd1)^~(4'd13)):((5'sd4)^(-3'sd2))));
  localparam signed [5:0] p5 = {{(3'sd0),(-5'sd7),(-5'sd7)},((2'd0)?(4'd6):(-3'sd1)),((6'd2 * (5'd10))&((2'd2)>=(2'd2)))};
  localparam [3:0] p6 = (-3'sd0);
  localparam [4:0] p7 = (((3'sd0)?(4'd1):(5'd5))%(2'd3));
  localparam [5:0] p8 = (|((+(((3'sd3)<(-4'sd4))&&((-4'sd6)&&(4'd3))))+((~(3'sd2))!=(-(4'd3)))));
  localparam signed [3:0] p9 = (({(4'sd2)}?{(-2'sd1),(3'd7),(3'd7)}:((3'd2)>>>(-4'sd5)))^((~^(5'd25))?((4'sd5)!=(5'd17)):((3'sd3)?(5'sd15):(4'd5))));
  localparam signed [4:0] p10 = ((2'd0)?(3'sd2):(3'sd2));
  localparam signed [5:0] p11 = (5'd2 * ((2'd0)<<<(4'd2)));
  localparam [3:0] p12 = (((5'd13)?(5'd8):(5'd15))?(-(&(|(-4'sd3)))):{3{(4'd15)}});
  localparam [4:0] p13 = ((((3'd4)>(3'd1))>={(5'd24)})?(((2'd3)?(5'sd3):(-4'sd7))^((5'd20)?(5'sd9):(4'd0))):(((5'sd12)?(2'd0):(5'd8))?(~^(3'd6)):((2'd3)!=(3'd4))));
  localparam [5:0] p14 = ((4'd11)|(((-5'sd6)?(4'd13):(3'd2))?{(2'd2),(-4'sd7),(4'd13)}:(3'd2)));
  localparam signed [3:0] p15 = (~&((6'd2 * (3'd6))^((3'd1)-(4'sd6))));
  localparam signed [4:0] p16 = {((5'd2 * (4'd2))-((4'd14)+(4'sd2))),{((2'sd0)!==(2'sd1)),{(2'd3),(-2'sd1),(5'sd2)}},{(~|(3'd0)),((-5'sd7)|(2'd3))}};
  localparam signed [5:0] p17 = (((-4'sd0)<((5'd29)?(5'd7):(5'd8)))==(((5'sd13)-(2'sd0))?((3'd0)||(-5'sd13)):((3'sd2)/(-2'sd0))));

  assign y0 = {({(4'd2 * $unsigned((b1!==b2))),($unsigned({p6,a0,p0})&&(b2>=p11)),((b3>=a1)+(p5>a0))})};
  assign y1 = {2{{{p7,p9},(4'd3)}}};
  assign y2 = (a0?b2:b2);
  assign y3 = ((p8>>>p11)?(p9?p2:p15):(&{1{p13}}));
  assign y4 = (|((p5>=p13)?(p4?p5:p0):(3'd3)));
  assign y5 = {1{{4{{a4,b3,b2}}}}};
  assign y6 = {3{a4}};
  assign y7 = {4{{p0,p17,b0}}};
  assign y8 = (({4{b4}}<=(p13<=b1))&&{4{(5'd2 * p6)}});
  assign y9 = ($signed(((3'd4)!==(b3>=b1)))!=(^{4{b1}}));
  assign y10 = ((p7>p0)&&(-{3{b4}}));
  assign y11 = $signed((5'sd8));
  assign y12 = (({2{b5}}?{3{b5}}:(p15?a0:a0))?{4{a0}}:({4{a5}}?{2{a2}}:{2{b5}}));
  assign y13 = {4{(~^($unsigned(a5)&&(a1&&b0)))}};
  assign y14 = (+(a2-b4));
  assign y15 = (((6'd2 * a2)==(p11<<<b3))&(6'd2 * (p2+a0)));
  assign y16 = ({3{p13}}&(p14!=a2));
  assign y17 = ((6'd2 * (!(p0>>b1)))^(&(~|(&(a0==p1)))));
endmodule
