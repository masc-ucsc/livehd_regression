module expression_00346(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-5'sd0)-(3'sd2))<<<((-5'sd2)&(-2'sd1)))>=((+(3'd0))?(3'd1):((3'sd2)?(-5'sd10):(-2'sd1))));
  localparam [4:0] p1 = (~|(((3'd5)?(3'd6):(5'd17))?((5'd25)?(3'd6):(5'd14)):(~&(4'd12))));
  localparam [5:0] p2 = (&((^(3'sd3))===((3'd7)+(3'sd0))));
  localparam signed [3:0] p3 = {1{(|{1{{4{(5'sd4)}}}})}};
  localparam signed [4:0] p4 = (-5'sd2);
  localparam signed [5:0] p5 = ({3{((3'd7)?(2'd3):(5'd13))}}?(^(~^((-3'sd3)?(-3'sd1):(4'd13)))):(((4'd5)?(3'sd2):(-4'sd7))?(&(5'd5)):((2'd2)?(2'd2):(2'd1))));
  localparam [3:0] p6 = {2{{3{((-2'sd0)!=(-5'sd11))}}}};
  localparam [4:0] p7 = {{4{(4'd7)}},{(2'sd1),(4'd7),(4'd3)},{(5'd4),(-2'sd0),(4'd9)}};
  localparam [5:0] p8 = (!{{(4'sd0),(3'd0)},(+(~&(-2'sd0))),{{(2'd2),(5'sd1),(-5'sd0)}}});
  localparam signed [3:0] p9 = (2'd3);
  localparam signed [4:0] p10 = ((5'd25)^~((4'sd7)>>(-2'sd0)));
  localparam signed [5:0] p11 = (^{1{(((-4'sd1)&(2'sd0))?((4'sd0)<(2'd3)):(&((-2'sd1)-(5'd28))))}});
  localparam [3:0] p12 = ((-(-2'sd0))>>>(4'sd5));
  localparam [4:0] p13 = {({(3'sd3),(2'd2)}===(4'd1)),(((2'sd0)>=(5'd12))&&((5'd21)>=(2'd3)))};
  localparam [5:0] p14 = {{{4{(3'd0)}},((5'd23)>>>(4'sd6)),{4{(3'd0)}}},{2{{2{(-4'sd5)}}}},{(~|{4{(4'sd1)}})}};
  localparam signed [3:0] p15 = ((((4'd8)?(-4'sd2):(-2'sd0))?((2'sd0)&&(4'd2)):((4'sd7)<<(4'sd0)))||(!(((3'sd1)==(4'sd1))?(~&(5'd6)):((-5'sd13)?(2'd1):(3'd4)))));
  localparam signed [4:0] p16 = {1{(3'd5)}};
  localparam signed [5:0] p17 = ((-2'sd1)||(2'd0));

  assign y0 = ((p13?p4:p12)!=((p15?p12:p10)+(p5<<p8)));
  assign y1 = (~^{(4'sd1),{{4{b1}},(3'sd0),{p11}},(-3'sd0)});
  assign y2 = $signed({2{$unsigned((((b3?a4:a0))+{a2,a1,b4}))}});
  assign y3 = {1{(~&{4{(b4!==b3)}})}};
  assign y4 = (((a4?a4:b1)<<<{2{a0}})<(4'd6));
  assign y5 = (~^(~(p11?p9:b3)));
  assign y6 = ((b2?p3:p10)?(~|(p12>>>a5)):(-(!(~b0))));
  assign y7 = (((~|p2)^(p9|p8))^(+(4'd3)));
  assign y8 = {2{$signed((&{2{$unsigned(p12)}}))}};
  assign y9 = (4'sd2);
  assign y10 = (^((4'd2 * (p8<=p0))?{(p4^p9),$signed({p4})}:($unsigned((p5?p0:a4))>>{(-3'sd3)})));
  assign y11 = {3{((-4'sd3)?(p13|p12):(+p11))}};
  assign y12 = $signed((((a1==a0)&&$unsigned((a4)))?({2{a3}}^(a0&b3)):{4{(a2==a5)}}));
  assign y13 = (~|((a2>=b5)!==(4'sd0)));
  assign y14 = (^(a5?p9:p9));
  assign y15 = (((((b4<=a5)*(~a2)))!==(&(~|(b1>=a1))))>(((~b2)|$signed(a5))|((p8>>a2)&&(a3!==b1))));
  assign y16 = {$unsigned((~|((a4?a5:p5)?(b1<<<a4):(4'd0)))),((a2===a5)?(-(&b4)):(&(&b1)))};
  assign y17 = $unsigned({((b2!==a1)?(p9>=p3):(p5<<a1))});
endmodule
