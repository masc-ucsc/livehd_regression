module expression_00637(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~^((~|(|(5'sd9)))<<<((3'd7)<=(-5'sd1))))^(!(|(((2'sd0)<=(4'sd3))!=(~^(~^(5'sd15)))))));
  localparam [4:0] p1 = (({1{{4{(4'd14)}}}}<<<{2{(2'd2)}})^({(2'd0),(5'sd6)}?((3'sd3)!=(2'd1)):((3'd0)^~(5'd25))));
  localparam [5:0] p2 = ((4'd2 * (2'd3))!={(3'd7),(-2'sd1)});
  localparam signed [3:0] p3 = {3{((&(3'sd3))==((4'd15)<<<(-3'sd1)))}};
  localparam signed [4:0] p4 = ({1{((5'd16)?{(3'sd0),(5'd29),(2'd2)}:((2'd0)!==(2'd3)))}}!==(((2'sd0)?(5'd10):(3'd0))?((5'd17)?(-3'sd1):(-5'sd1)):{(2'd2),(5'd31),(-4'sd3)}));
  localparam signed [5:0] p5 = (((4'd10)^~(-2'sd0))>>{{2{(-2'sd0)}}});
  localparam [3:0] p6 = {(!(~(~|((2'sd1)||(2'd0)))))};
  localparam [4:0] p7 = (-5'sd10);
  localparam [5:0] p8 = ((!({3{(-3'sd1)}}-((5'd5)>(5'd16))))<<(-5'sd10));
  localparam signed [3:0] p9 = ({2{{4{(5'd21)}}}}>=({(4'sd6),(2'd0)}&(&(2'd0))));
  localparam signed [4:0] p10 = {{2{{1{(-2'sd1)}}}},(|{(5'd30),(2'd1),(2'd1)}),(~&{4{(2'sd1)}})};
  localparam signed [5:0] p11 = {{((2'sd1)||(-2'sd1)),((-3'sd1)<<(3'sd3)),{3{(5'd19)}}},((4'd2 * (5'd9))<((-4'sd7)>(-3'sd3)))};
  localparam [3:0] p12 = ((-5'sd6)<<(2'd0));
  localparam [4:0] p13 = (3'd1);
  localparam [5:0] p14 = ((&((4'd6)>=(-2'sd0)))%(4'd7));
  localparam signed [3:0] p15 = {(4'd12),(-5'sd4),(2'sd0)};
  localparam signed [4:0] p16 = (-5'sd6);
  localparam signed [5:0] p17 = (5'd25);

  assign y0 = $signed((a2?b1:a1));
  assign y1 = (5'sd13);
  assign y2 = $unsigned(((b2?a3:b2)&&$signed(a2)));
  assign y3 = ((+(p10||a4)));
  assign y4 = (|(+{{(~{b1,p5})},(4'sd4),(^(~&(-5'sd9)))}));
  assign y5 = (-$signed(((3'd4)?(3'd6):(2'd0))));
  assign y6 = ((-5'sd4)^~(4'd12));
  assign y7 = (($unsigned({{b2,b2,a4},(~&b0),(b4?a1:a0)}))&$signed(({{a1,b3},$signed(a4)}==(~|(4'd2 * b0)))));
  assign y8 = (~&(&((+(+(+(-(|(~(~&p7)))))))>>>(|((~|(^a5))^~(-(b0||a1)))))));
  assign y9 = {(~&{(p0<a5),(a2<<p16)}),(&{(a1>>p0),(+(&b0))})};
  assign y10 = (-4'sd2);
  assign y11 = $unsigned($signed((+(+(^(-5'sd0))))));
  assign y12 = {{4{(+a5)}},{4{{1{p11}}}},$unsigned(((b0==a3)<=(p11<<<p9)))};
  assign y13 = ((2'd2)>=(a0?p0:a2));
  assign y14 = (-{(&p0),(p1<p17),{p6,a5}});
  assign y15 = ((~&(((a3<a3)&&(-2'sd1))>(4'd12)))===(~(&((a2<=a4)*(a5*a5)))));
  assign y16 = (((b2&a2)!==((b4>=b0)))===(((~^b0)|(b0<=a2))));
  assign y17 = (~^(~(a1^b2)));
endmodule
