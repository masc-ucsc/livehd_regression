module expression_00872(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((4'd10)!==(4'd1)),((-4'sd7)?(2'd1):(2'sd0))};
  localparam [4:0] p1 = (^(4'sd7));
  localparam [5:0] p2 = ((3'd4)?(2'd3):(5'd24));
  localparam signed [3:0] p3 = ((2'sd1)==(-4'sd3));
  localparam signed [4:0] p4 = (-5'sd4);
  localparam signed [5:0] p5 = {(((4'd14)||(2'sd0))?((5'sd6)?(2'sd0):(-3'sd0)):(6'd2 * (4'd4))),(((3'd7)>>>(3'sd1))&{(5'd7),(2'd3)})};
  localparam [3:0] p6 = {3{(5'sd10)}};
  localparam [4:0] p7 = (^((^((2'sd0)&(2'd1)))<<{(4'd13),(4'd6),(2'd0)}));
  localparam [5:0] p8 = (~{((5'd2)?(2'sd0):(4'd7)),(~&(4'd13)),((3'd6)?(4'sd7):(-2'sd1))});
  localparam signed [3:0] p9 = (~|((+((-5'sd6)<<<(5'd23)))?(|((2'd1)===(4'sd6))):((4'd2)?(5'd19):(5'sd11))));
  localparam signed [4:0] p10 = (|(|{3{(&(~|((5'sd7)?(-5'sd2):(3'sd3))))}}));
  localparam signed [5:0] p11 = (&(!(~|(&(3'd3)))));
  localparam [3:0] p12 = {{{{{(-4'sd5),(5'sd9),(2'd3)},{(2'sd1)},{(4'sd3)}}},{{{(2'sd0)},{(5'd23)},{(4'd15)}}}}};
  localparam [4:0] p13 = (-4'sd6);
  localparam [5:0] p14 = ({4{(2'sd0)}}^~(5'sd2));
  localparam signed [3:0] p15 = (!(^{3{(~^(-5'sd13))}}));
  localparam signed [4:0] p16 = (~|{((~|(5'd6))-((2'd3)>(3'd4))),(~&((-5'sd14)>=(2'd0)))});
  localparam signed [5:0] p17 = (~^((((-3'sd1)?(-2'sd1):(2'sd1))!={(3'd3),(-4'sd5),(2'd3)})|(&(~&((-5'sd12)===(-3'sd0))))));

  assign y0 = (b2||b0);
  assign y1 = {p15};
  assign y2 = ({1{(4'd14)}}?$unsigned((p17?p2:p16)):(5'sd6));
  assign y3 = (~&(-(2'd3)));
  assign y4 = $signed({$signed((4'sd4)),(!(~&$signed({a3,a1,b2}))),(~&(~{b3,a2}))});
  assign y5 = (&{(6'd2 * (b0?a0:b1)),{1{(a1>>p1)}},((b1^p12)==(|b1))});
  assign y6 = ((((b3+b2)!==(b1+b1))>>>(p0?p3:p8))<((+(&(a3?a2:a2)))>>>((p6/p11)>>(p4?p16:p13))));
  assign y7 = (({p6,a0,p5}<=(|(a0!==b5)))<((a2!==b1)>{p17,a3,p1}));
  assign y8 = (&(~&{3{(~|{p5,p16,p15})}}));
  assign y9 = (~{(((a3>=b3)?{a3,a4}:(b4>a4))!=((b2?p11:p5)^(4'sd2)))});
  assign y10 = {(^(^{a4,p17,p12})),$unsigned((&(~|b2))),{(p17&&b2),(a1)}};
  assign y11 = (~|({(!(-4'sd3)),(-2'sd1)}?{1{(~^(~^(-4'sd5)))}}:(-({1{a3}}?(~&a0):(~&a2)))));
  assign y12 = (|((!(~&((~|p17)>>>(p5||p5))))<<{4{{1{p7}}}}));
  assign y13 = (~&(-(~&p1)));
  assign y14 = ((((p4<p1)<<<(p0^~p11))-($signed((a1+b2))===$signed((a4<b1)))));
  assign y15 = (-2'sd0);
  assign y16 = (((b5?a4:b3)?(b0<<a2):(a0?b2:b1))===((-((b0>=a0)^(b3?b2:a4)))!==({a1,b2}<<(a5-a0))));
  assign y17 = {(~^(!{a3,a4,b1}))};
endmodule
