module expression_00825(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^((((-5'sd3)||(-3'sd1))-{4{(4'd5)}})==(((3'd5)&(3'd5))!==(-2'sd1))));
  localparam [4:0] p1 = {4{(((3'd4)>(4'd14))>>>((2'sd1)==(3'd6)))}};
  localparam [5:0] p2 = (5'd10);
  localparam signed [3:0] p3 = ((((3'sd1)<=(3'sd3))<((3'sd0)-(2'd1)))>>{(4'd13),(2'sd0),(5'd13)});
  localparam signed [4:0] p4 = (4'sd3);
  localparam signed [5:0] p5 = {1{{1{{((4'd13)>(-2'sd0)),((-4'sd5)&&(5'd31)),(~&(2'd3))}}}}};
  localparam [3:0] p6 = (4'd2 * ((5'd15)<<(4'd2)));
  localparam [4:0] p7 = (({((2'd0)!==(4'd13)),{(2'd0),(5'sd15)}}<{(5'd2 * (4'd5)),((4'd14)<=(-4'sd4))})<(-3'sd3));
  localparam [5:0] p8 = {4{(5'sd0)}};
  localparam signed [3:0] p9 = (({1{(3'd1)}}?{2{(3'd6)}}:((3'd3)<<(-4'sd0)))>=((5'd28)===((3'sd2)?(4'sd2):(4'd11))));
  localparam signed [4:0] p10 = (^(~^(~(^(~&(-(-2'sd0)))))));
  localparam signed [5:0] p11 = ({(4'd2 * (4'd4)),((-4'sd2)>>(-2'sd0)),{(5'd3)}}<=(4'd2 * ((4'd14)||(3'd3))));
  localparam [3:0] p12 = (5'd0);
  localparam [4:0] p13 = {((3'd2)?(5'd23):(4'd3)),((-5'sd14)>>(-2'sd0)),((3'd7)&(5'sd13))};
  localparam [5:0] p14 = (({2{(5'sd12)}}&(+(5'd2 * (5'd2))))||{2{{1{((4'sd0)===(-4'sd0))}}}});
  localparam signed [3:0] p15 = (|(&(4'd15)));
  localparam signed [4:0] p16 = {1{(~&(3'sd3))}};
  localparam signed [5:0] p17 = (~{1{{4{(~|{4{(-5'sd14)}})}}}});

  assign y0 = (((!a1)-(3'd4))!==(4'd8));
  assign y1 = (3'd4);
  assign y2 = (((5'd3)%b5)&((6'd2 * p0)*(p12!=p8)));
  assign y3 = {{1{(!(b3>>b0))}},{{a0,b0,p15}},(2'd1)};
  assign y4 = (-5'sd1);
  assign y5 = (5'd9);
  assign y6 = ({1{p3}}?(~|a1):(+a2));
  assign y7 = (^{3{p7}});
  assign y8 = ((+(^{2{{2{(^$signed((~&p6)))}}}})));
  assign y9 = ((a2?b1:b3)>=(p12?b2:b3));
  assign y10 = {3{({2{p7}}>>>(a2===a4))}};
  assign y11 = (((b2-b5)|(-a2))>>>$signed($signed((b5!==a5))));
  assign y12 = (~|{4{{4{p9}}}});
  assign y13 = (((p14/p4)>=(b1<=a1))+((p3>>>p12)&(5'd2 * p2)));
  assign y14 = {2{(5'd31)}};
  assign y15 = (-((|(&{4{a3}}))<<<(+(~&{1{a2}}))));
  assign y16 = (~^((~(({p9,p4,p7}^(p0<<b3))!=((~p10)<<(-p12))))^(3'd0)));
  assign y17 = (+{(b0?p5:b0)});
endmodule
