module expression_00012(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(3'd4),(2'd2),(5'd15)}!==((3'd0)&&(2'd3)));
  localparam [4:0] p1 = {1{({{(2'sd1),(5'd3),(4'd15)}}?(((-2'sd1)>(-3'sd3))^~((2'd2)>>(-2'sd1))):({(5'd10),(4'd7)}-{(-5'sd6),(2'd2),(3'd7)}))}};
  localparam [5:0] p2 = ((4'd1)?(3'd2):(4'd1));
  localparam signed [3:0] p3 = ((((-2'sd0)-(2'd2))^(|(5'd18)))-(6'd2 * (+((2'd0)^~(5'd25)))));
  localparam signed [4:0] p4 = (3'd3);
  localparam signed [5:0] p5 = (3'd0);
  localparam [3:0] p6 = {1{(((4'd1)<<<(4'd12))>>>{1{(4'd8)}})}};
  localparam [4:0] p7 = (((3'd6)?(3'd2):(4'd2))?(4'd7):(-4'sd6));
  localparam [5:0] p8 = (((4'd4)^(-4'sd6))<((3'd2)|(2'sd1)));
  localparam signed [3:0] p9 = ({(3'd1),(2'd0)}!=={(5'd23)});
  localparam signed [4:0] p10 = (~&((~^((2'sd0)==(4'd13)))?((4'sd1)<<(-2'sd1)):(~^(~|(-3'sd2)))));
  localparam signed [5:0] p11 = {4{(5'd2)}};
  localparam [3:0] p12 = ((3'd7)&&(-4'sd7));
  localparam [4:0] p13 = ((+(&((-3'sd1)<=(3'd7))))<<((~(-4'sd2))?((5'sd6)?(3'd7):(5'd16)):((5'sd5)?(3'd7):(5'd6))));
  localparam [5:0] p14 = (~|{1{({1{(&(-{2{(5'd31)}}))}}==(6'd2 * (+(!(5'd26)))))}});
  localparam signed [3:0] p15 = ((((2'd3)==(3'sd1))<((-5'sd3)===(4'd4)))<(~|(~((&(4'sd1))+((3'd4)>>>(-5'sd5))))));
  localparam signed [4:0] p16 = (2'sd0);
  localparam signed [5:0] p17 = ((((2'sd0)?(2'sd0):(-5'sd12))<=((5'd15)>(5'd14)))>>(-3'sd1));

  assign y0 = {{(-5'sd5),{(3'd6)}},(-5'sd5)};
  assign y1 = {{2{(~|(&p3))}},({{4{p14}}}),(~|$unsigned({1{(3'sd1)}}))};
  assign y2 = ({((-5'sd1)&{p11}),(-3'sd1)}=={(b5>=p11),(b1==p17),(p1-p6)});
  assign y3 = (p4?p10:a3);
  assign y4 = (~&((((^b0)>=(|a2))+(2'sd1))!=(~|((4'sd5)<<<{4{b0}}))));
  assign y5 = (((a1?p10:b0)?(5'd11):(-3'sd3))?(($signed((a5?a1:a5)))):$signed($unsigned((a5?b2:a4))));
  assign y6 = {2{({{p11,p14,p2},(p9&p0),(~^p11)}>>{((p17&&p0)!={1{p16}})})}};
  assign y7 = {1{(((p13-p11)!=(p0?b1:p12))^~((p17&&b1)>={1{a3}}))}};
  assign y8 = (-2'sd0);
  assign y9 = $unsigned($signed((5'd23)));
  assign y10 = (-((a1?p8:b3)?{p9,b4}:(p17?p12:p16)));
  assign y11 = (~&{2{b4}});
  assign y12 = (!((4'd2)^~(4'd12)));
  assign y13 = $unsigned($unsigned((b0&a2)));
  assign y14 = (((a5|b0)?{2{p14}}:$unsigned(a4))<<($signed(b1)>>(a5&b0)));
  assign y15 = (&(b2<=p6));
  assign y16 = ({p5,p10}-(p1<b4));
  assign y17 = (^{{{p9},(|p7),(~p17)},(~&{{{p16,p7,p15}}}),(&((~^p14)<<(p0>>>p11)))});
endmodule
