module expression_00662(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~^((4'd12)===(3'd4)))>=((3'd2)===(-4'sd5)))>={(&({(4'd8),(4'd5)}>=(|(5'd17))))});
  localparam [4:0] p1 = (&{(^(5'd9)),(+(3'sd3)),{(3'sd3),(4'd4),(-2'sd0)}});
  localparam [5:0] p2 = {(3'sd2)};
  localparam signed [3:0] p3 = (-3'sd0);
  localparam signed [4:0] p4 = ((!(-(3'd7)))>={((2'd1)>>(4'd5))});
  localparam signed [5:0] p5 = {(~|(~^(~^(~(5'd16))))),{{(-2'sd0),(5'd3)},(|(-2'sd0))},(~&{{(-3'sd1),(-5'sd4)},(~(3'sd0))})};
  localparam [3:0] p6 = {{{2{(5'd6)}}},(~&(!((4'd0)==(3'd3)))),{4{(2'd1)}}};
  localparam [4:0] p7 = ((-4'sd3)?(2'd2):(3'sd2));
  localparam [5:0] p8 = ((^(3'd3))!=(~^(4'd9)));
  localparam signed [3:0] p9 = ((+(((5'sd9)==(5'sd7))<<<((4'sd6)|(2'sd1))))<<(((2'sd0)<=(-2'sd0))<<(^(3'd6))));
  localparam signed [4:0] p10 = ((-4'sd2)!==(2'sd1));
  localparam signed [5:0] p11 = (((2'sd1)<(-4'sd7))?{(3'd6),(2'd3)}:((2'sd1)&&(5'd24)));
  localparam [3:0] p12 = {(^(-((5'd27)|(2'd2)))),{2{((2'd3)||(-4'sd2))}},(3'sd2)};
  localparam [4:0] p13 = (5'd20);
  localparam [5:0] p14 = ((-3'sd2)<{(((-2'sd1)!==(5'd8))||{(-3'sd3)})});
  localparam signed [3:0] p15 = ((4'd7)===(-4'sd2));
  localparam signed [4:0] p16 = (-5'sd15);
  localparam signed [5:0] p17 = ((4'd2 * ((2'd3)*(5'd14)))==(((4'sd7)?(2'sd1):(5'd5))?((-5'sd0)<<<(-3'sd3)):((-4'sd2)==(4'sd2))));

  assign y0 = (&(-3'sd0));
  assign y1 = (4'd12);
  assign y2 = {1{({4{{1{a5}}}}!==((^(b3<<b4))-(&{2{a2}})))}};
  assign y3 = ((3'd1)===(b1|a2));
  assign y4 = ((((~((&(-$signed(p11)))>={4{a3}}))<((~^(~^{3{{3{p6}}}}))))));
  assign y5 = {p9,a2,p0};
  assign y6 = {({4{b1}}?(a3?b1:b5):{b4,a3,b4})};
  assign y7 = (~&(((-(a4?a0:b1))?(+(b5?b5:a4)):(+(~b4)))<<((~^(b5==a2))?(|$signed(a5)):(a2?a4:a0))));
  assign y8 = ((a4%p14)/a0);
  assign y9 = (^{1{$unsigned((&(!(~|{(~&{3{p13}}),{4{p7}},{3{(b5>p16)}}}))))}});
  assign y10 = $unsigned((4'd8));
  assign y11 = (^(({a4,b5,a4}<<({p4,b0,p13}|(3'sd0)))&&(!(+((p7-b3)==(2'd0))))));
  assign y12 = ((p0?p12:a1)<{(a2?p16:p4)});
  assign y13 = ({1{(p7?p1:p16)}}<={2{p15}});
  assign y14 = (^((+(&(^(~&(a0!=b3)))))<=(^(^{(-(^b1))}))));
  assign y15 = (5'd2 * {3{p2}});
  assign y16 = (|((p12>>p17)!=(&(+p17))));
  assign y17 = {((4'sd3)||(b2?a2:a5))};
endmodule
