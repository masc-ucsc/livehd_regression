module expression_00718(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^{3{(!((4'sd1)-(3'd6)))}});
  localparam [4:0] p1 = (((~|((5'sd14)&&(5'd19)))^(+(-4'sd7)))<=(|(((-3'sd0)!==(5'sd15))|((3'sd1)===(3'd6)))));
  localparam [5:0] p2 = (3'd2);
  localparam signed [3:0] p3 = (+((&(5'd2))===((~|(|(2'sd0)))^(-((5'd23)^(2'd1))))));
  localparam signed [4:0] p4 = (~^(~|(^(~|(~|{(4'd9),(-2'sd1)})))));
  localparam signed [5:0] p5 = (5'd1);
  localparam [3:0] p6 = {((5'd15)<<<(2'd1)),((5'sd6)-(2'sd1))};
  localparam [4:0] p7 = {(2'd0)};
  localparam [5:0] p8 = (^(((-3'sd2)<<(2'd0))^((-5'sd15)^~(4'sd1))));
  localparam signed [3:0] p9 = (({4{(3'd2)}}>=(4'sd7))<=(-2'sd0));
  localparam signed [4:0] p10 = ({4{(2'sd1)}}|((4'd13)^~(5'sd14)));
  localparam signed [5:0] p11 = {(5'sd1)};
  localparam [3:0] p12 = (~&(({(3'd0),(3'd2),(4'sd5)}==(^(2'd2)))<(+(~(4'd2 * (5'd1))))));
  localparam [4:0] p13 = {1{(((2'sd0)>>>(2'sd1))&{((-4'sd3)||(-2'sd1))})}};
  localparam [5:0] p14 = (((4'sd7)==(-3'sd0))+(5'd2));
  localparam signed [3:0] p15 = {3{{2{{(3'sd2),(5'd14),(3'd4)}}}}};
  localparam signed [4:0] p16 = (((2'd2)?(-5'sd12):(3'd3))?(~&{1{(5'd5)}}):{2{(2'sd1)}});
  localparam signed [5:0] p17 = ((((5'sd10)+(-4'sd5))&&{1{((2'd3)==(-2'sd0))}})>=((4'd2 * (2'd3))=={4{(2'd3)}}));

  assign y0 = {2{a4}};
  assign y1 = {(^(+{b5})),{{a2,p17}}};
  assign y2 = ((b2>>a2)===(3'sd3));
  assign y3 = ((5'sd6)<=(((4'd12)=={3{p9}})+({1{p16}}|(a2===b3))));
  assign y4 = (-4'sd0);
  assign y5 = (p10?b2:p10);
  assign y6 = {({4{p4}}|{a0,p9})};
  assign y7 = {{(~(~^a0))}};
  assign y8 = (|((5'd22)?((p8?p13:p12)&(p9?a2:p16)):({4{p13}}^(-3'sd3))));
  assign y9 = ({$unsigned({{b4},(~|p14)}),{4{b3}}});
  assign y10 = (4'd3);
  assign y11 = (-4'sd2);
  assign y12 = ((~^{3{{3{b1}}}})===({$unsigned(a3),(a3&&b3)}-(~^(~^{4{b1}}))));
  assign y13 = {4{a2}};
  assign y14 = ((~^{((b4<<<b4)|(b2|b0))})<<((-(~{a1}))-(^{a3,p10,p11})));
  assign y15 = (((a1?a5:a0)?{1{{4{b0}}}}:{1{(b0?a1:a4)}})<<($signed((b4))?$unsigned((a4?b2:a5)):(p3-b2)));
  assign y16 = (($signed(p5)?{4{a0}}:{p13})|((a1?p15:p6)?(a4==p4):(b0&&a0)));
  assign y17 = (&(6'd2 * $unsigned((!b2))));
endmodule
