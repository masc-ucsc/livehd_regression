module expression_00916(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{{1{((3'sd1)==(-4'sd5))}}}};
  localparam [4:0] p1 = {4{(3'd7)}};
  localparam [5:0] p2 = (4'sd4);
  localparam signed [3:0] p3 = ((5'd26)?(5'd7):(4'd9));
  localparam signed [4:0] p4 = (^(&(-2'sd0)));
  localparam signed [5:0] p5 = ({2{(5'sd15)}}==(-3'sd2));
  localparam [3:0] p6 = ({(~(~|(4'd6))),((4'd1)>>>(-3'sd2))}<={2{{(-2'sd1),(2'sd1)}}});
  localparam [4:0] p7 = {(((&(5'd15))>((-2'sd1)?(5'sd8):(4'd15)))>(~|((-3'sd3)?(3'd0):(-2'sd1))))};
  localparam [5:0] p8 = {1{(&(((-2'sd1)^~(3'd7))&&((4'sd7)-(-2'sd1))))}};
  localparam signed [3:0] p9 = (3'sd1);
  localparam signed [4:0] p10 = ((!(4'd12))?(&(-3'sd3)):(4'd2 * (5'd28)));
  localparam signed [5:0] p11 = ((5'd21)?(-2'sd1):(2'd2));
  localparam [3:0] p12 = (((((4'd12)&(3'sd0))/(2'd3))|(((4'sd3)&(-3'sd2))>>>((-2'sd1)%(4'd3))))>>>(((5'd3)&(5'd18))%(-3'sd2)));
  localparam [4:0] p13 = ((((4'd13)>>(4'd8))!=(-4'sd7))-((-(3'd2))^~((5'd10)===(-4'sd6))));
  localparam [5:0] p14 = ({2{(4'd14)}}<((3'd2)&(-2'sd0)));
  localparam signed [3:0] p15 = (+(!(^(~^(~&(!(^(~&(|(~^(~&(&(5'd11)))))))))))));
  localparam signed [4:0] p16 = ((3'd1)?(^(-3'sd0)):((4'sd0)?(-5'sd7):(-4'sd6)));
  localparam signed [5:0] p17 = (2'sd1);

  assign y0 = (|$signed(((!((4'sd1)?$signed($signed(p17)):(p4^p6)))-((^(a4?a2:b5))^~$unsigned((b4?p15:p9))))));
  assign y1 = ({(-3'sd0),{4{b3}},{3{a5}}}?{(a3?b5:b0),{b2},{4{a4}}}:{{1{(5'd13)}}});
  assign y2 = ((a5>b0)&&(a1!=p2));
  assign y3 = (((b3^~b4)==(a3?b1:b1))>((b0?b2:a5)&{a5,b3}));
  assign y4 = (b5?a2:b0);
  assign y5 = ($unsigned(p12)<<(+p10));
  assign y6 = (b3&b0);
  assign y7 = (!$unsigned({p15}));
  assign y8 = (a1>>b3);
  assign y9 = {1{(&((!{4{p8}})?((&p16)?(b0+b0):{p2}):(+((a4>=p6)==(~a4)))))}};
  assign y10 = ((~|(p9<<a0))?(a2*a4):(|(p0%b3)));
  assign y11 = {4{({p12,p10}!=(p8<<<a5))}};
  assign y12 = (~$unsigned((((~|(a4&a1))^~{a5,b5,b0}))));
  assign y13 = ((2'sd0)<=(-2'sd0));
  assign y14 = (~|p0);
  assign y15 = ($signed(a5)*$unsigned(a3));
  assign y16 = {{(p4<a1)},(p13?a1:p6),(a4==a5)};
  assign y17 = {{($unsigned({a5})?(+(^b4)):{b1,p0,p10}),(-{(p4>a4),{p15},{p15}})}};
endmodule
