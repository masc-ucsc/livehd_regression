module expression_00934(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd3);
  localparam [4:0] p1 = (|(((~(-3'sd1))!=((5'd24)?(5'd31):(3'd7)))>>>((2'sd0)?(2'd2):(3'd0))));
  localparam [5:0] p2 = (4'd8);
  localparam signed [3:0] p3 = (-2'sd1);
  localparam signed [4:0] p4 = ((((2'd3)>>>(2'sd1))%(4'sd1))||(((2'd3)>=(-4'sd5))+((5'd20)==(-5'sd1))));
  localparam signed [5:0] p5 = ({2{((5'd18)<=(4'd0))}}>>((-3'sd0)+{(4'd5)}));
  localparam [3:0] p6 = ((((4'd10)<(5'd7))^~((-5'sd1)>>>(-3'sd0)))+(((4'sd0)||(2'sd0))|((3'sd0)^(5'd19))));
  localparam [4:0] p7 = ((~^(+{3{(-5'sd6)}}))>{2{((3'd1)!==(-2'sd1))}});
  localparam [5:0] p8 = (-3'sd2);
  localparam signed [3:0] p9 = (~|(|{((3'd1)?(5'd0):(2'd3)),((2'sd1)+(5'sd9)),(~(!(3'sd3)))}));
  localparam signed [4:0] p10 = (({4{(5'sd15)}}?((4'sd2)?(4'd5):(2'sd1)):(~(2'd2)))-(((4'sd4)?(3'sd0):(5'd22))|{3{(-3'sd2)}}));
  localparam signed [5:0] p11 = ((!(4'd0))>>((5'sd7)|(-2'sd0)));
  localparam [3:0] p12 = ((4'sd1)<={3{(-4'sd7)}});
  localparam [4:0] p13 = (({(4'd13),(-2'sd0),(3'd3)}^~{4{(2'sd1)}})||({3{(3'd5)}}<=((-4'sd2)+(2'd1))));
  localparam [5:0] p14 = {({(3'd4),(4'sd7)}<<<((3'd5)&(4'sd6))),{{(2'd2),(3'sd3)},((2'sd0)===(5'd22))}};
  localparam signed [3:0] p15 = (5'd14);
  localparam signed [4:0] p16 = {(-((5'd23)&&((4'sd1)<=(4'd11)))),(2'd0),(~&({(4'd6)}!=(|(2'sd0))))};
  localparam signed [5:0] p17 = ({(((-5'sd9)+(3'd4))^~(!(-2'sd1)))}+({(3'd6)}<((-5'sd10)?(5'd17):(5'sd3))));

  assign y0 = (((2'd1)==(5'd4))<<<((~(~|p6))*(!(p16%p1))));
  assign y1 = (!(a3&b2));
  assign y2 = (~|(((a1?a1:b5)*(b2>>>a3))?(-(3'sd3)):((3'sd1)-(3'sd1))));
  assign y3 = ((~^(~|a3))?(a2<b1):(~(b0==a2)));
  assign y4 = (4'sd7);
  assign y5 = {3{(~|(~&((p6<<p7)?(p2?a2:p8):(&b3))))}};
  assign y6 = (^(~{((!(p16+p15))|(~&(a1|p13))),(((p1!=a2)>(a3<p17))>$signed((^(~p14))))}));
  assign y7 = (~((&$signed(p6))));
  assign y8 = {2{(3'd7)}};
  assign y9 = (~^(&$unsigned((~(-$unsigned((~|($unsigned(((a3-b3)))===((b4>>>a3))))))))));
  assign y10 = ((^((~(~p17))<<(~&{b1,p15})))>>(!(~((b2<=a3)+(p10+p8)))));
  assign y11 = {({1{a4}}?{4{a2}}:$unsigned(a1))};
  assign y12 = ($signed($signed({2{p6}}))<((p5?a4:a0)!=(-5'sd6)));
  assign y13 = ((((p16?a2:b1)?{p11,b5}:(a2!==b5))!=((b5)&(~&p5)))<<<(6'd2 * (a1<<p8)));
  assign y14 = ((({2{b1}}!==$signed(a2))===($signed(a0)|(a4===b2)))<(({1{b2}}?(b2?a4:p7):$unsigned(b1))<<<{3{(b5?b2:p8)}}));
  assign y15 = (({4{b1}}&((+b4)+{2{b2}}))<<<((~(|{2{a1}}))===((a5===b2)>>>{1{a5}})));
  assign y16 = (&(!(|{1{p17}})));
  assign y17 = ((((b5?b4:b3)&(b2?p15:a0))<<{3{b1}})<(((a4?a1:p8)<(p1?p2:b1))!=(p7?a1:a3)));
endmodule
