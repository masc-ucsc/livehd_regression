module expression_00759(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^(((2'd2)?(5'd30):(3'sd1))?((2'sd0)?(2'sd1):(4'sd6)):((4'sd5)?(2'sd1):(4'd6))));
  localparam [4:0] p1 = (+{3{(^{(2'd0),(-5'sd15),(2'd2)})}});
  localparam [5:0] p2 = ({((5'd18)&&(2'sd1)),{(-4'sd2),(2'sd1)},{(3'sd1),(4'd14),(2'd0)}}<{3{((4'sd5)!==(2'sd1))}});
  localparam signed [3:0] p3 = (~^(~|{3{((-2'sd0)>(3'd0))}}));
  localparam signed [4:0] p4 = ((4'd1)&{4{(2'd1)}});
  localparam signed [5:0] p5 = ({((-3'sd3)==(5'd3)),(-4'sd2)}>>(((4'd12)!=(3'd6))===((4'd2)^(-2'sd1))));
  localparam [3:0] p6 = {4{{(3'd7),(-4'sd3),(5'sd4)}}};
  localparam [4:0] p7 = (|{{((-4'sd1)?(5'd9):(2'd0)),((2'd3)?(2'd3):(4'd4))}});
  localparam [5:0] p8 = {1{{2{(3'd3)}}}};
  localparam signed [3:0] p9 = {((3'd7)?(5'sd14):(-2'sd1)),{(3'd0),(5'd25),(5'sd0)}};
  localparam signed [4:0] p10 = (-(-(-{{(3'd7),(3'd6),(-5'sd2)},(~((5'sd5)?(4'sd1):(4'sd6))),{((-4'sd0)?(2'd0):(-5'sd15))}})));
  localparam signed [5:0] p11 = {(((3'd3)^~(4'sd5))^~{4{(-5'sd13)}}),((!(2'd1))+{(4'd0),(4'd15),(-4'sd5)})};
  localparam [3:0] p12 = ((((2'sd1)>(4'd14))|(^(!(5'sd5))))>((-((2'sd1)?(4'd7):(5'sd10)))<={(-4'sd3),(5'sd6)}));
  localparam [4:0] p13 = (4'd5);
  localparam [5:0] p14 = ({{(3'sd2),(-4'sd6)}}!=(((-4'sd5)>=(5'sd0))>>((4'd2)<<<(2'd0))));
  localparam signed [3:0] p15 = ((-4'sd2)?(5'd15):((4'd3)?(-4'sd6):(3'd4)));
  localparam signed [4:0] p16 = (^(4'd2 * {(3'd2),(3'd3),(5'd23)}));
  localparam signed [5:0] p17 = {(~&(((5'd30)-(4'd15))>>>{(5'sd3),(-4'sd5),(2'd3)})),{{(4'sd0)},{(3'd1),(5'd26)},((-2'sd0)||(2'sd1))}};

  assign y0 = {4{a4}};
  assign y1 = {(4'd2 * (b0>>a1)),{{(a2>>b4),(!b3)}}};
  assign y2 = {2{{1{{4{{1{p11}}}}}}}};
  assign y3 = (4'sd5);
  assign y4 = ((a4+b4)?(a5&&b4):(b2&&b0));
  assign y5 = (((p10!=p17)>>>(p8&b0))^((p15*p3)+(a2*p1)));
  assign y6 = {2{{1{(a3?a0:p3)}}}};
  assign y7 = ($unsigned((-3'sd1))>((5'd2 * p12)/b0));
  assign y8 = (~&{{3{{2{(p4?a4:p6)}}}}});
  assign y9 = $unsigned(((3'd0)|(-4'sd6)));
  assign y10 = ({1{a4}}==(+p16));
  assign y11 = $signed({(({2{a0}})>>>{1{{p2,a5}}})});
  assign y12 = (((a2?a2:p12)||(p13>>>p13))&&{3{{3{a0}}}});
  assign y13 = ($unsigned($unsigned({4{a0}}))==((p13==a1)));
  assign y14 = ((!(6'd2 * a2))-(5'd2 * a1));
  assign y15 = ($unsigned({{{3{{a2,p13,p8}}}},{(p17),$signed(a4),(a0===a2)}}));
  assign y16 = ({3{(6'd2 * b2)}});
  assign y17 = ($unsigned((4'd13))?$signed((b5?b0:b5)):{4{b2}});
endmodule
