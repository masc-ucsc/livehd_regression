module expression_00678(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{({1{(((5'd5)&(-2'sd0))||((3'd5)|(5'd28)))}}>(4'd4))}};
  localparam [4:0] p1 = (({(4'd1),(3'd4)}||((3'sd2)<=(-2'sd1)))&{({(3'd7),(5'sd15),(2'd2)}?((-2'sd0)|(2'sd1)):((5'd20)?(2'd2):(2'sd0)))});
  localparam [5:0] p2 = {2{{{(4'd5),(5'sd0)},(3'd2)}}};
  localparam signed [3:0] p3 = (+((^(((-5'sd7)===(-3'sd0))===((3'd7)|(-4'sd5))))===(((3'sd2)+(3'd7))<((4'd2)>>(-5'sd15)))));
  localparam signed [4:0] p4 = (~|(-4'sd0));
  localparam signed [5:0] p5 = (-3'sd2);
  localparam [3:0] p6 = (3'sd1);
  localparam [4:0] p7 = (^{3{{3{(4'sd5)}}}});
  localparam [5:0] p8 = {4{{2{(4'd2)}}}};
  localparam signed [3:0] p9 = (({2{(3'sd1)}}<=((-4'sd1)^(5'sd10)))<<(((-4'sd2)>(4'sd1))>((4'd9)>(2'sd0))));
  localparam signed [4:0] p10 = (((4'sd1)?(5'd14):(3'd6))<<(~^((5'd17)>>(3'd7))));
  localparam signed [5:0] p11 = ({(-5'sd15),(2'sd1)}>=(5'd21));
  localparam [3:0] p12 = (!(-3'sd2));
  localparam [4:0] p13 = {(~&{(-4'sd7),(-3'sd1),(2'd2)}),({(4'd0),(-4'sd2),(2'd2)}&&((2'd2)?(5'd20):(5'd29))),((2'sd0)?(4'sd5):(2'd0))};
  localparam [5:0] p14 = {(((~|(3'd1))?((2'sd0)>(2'd2)):((-5'sd14)?(4'd3):(4'd13)))||(+((&(2'd1))+((-4'sd4)|(4'd11)))))};
  localparam signed [3:0] p15 = (((4'd2 * ((4'd10)+(4'd9)))<=(((3'd1)+(-4'sd0))^~((5'd15)==(-3'sd2))))>>>((((-4'sd4)!==(4'd8))>>>((-2'sd0)+(3'd7)))<<<(((-2'sd1)&&(2'd3))<<((3'sd3)>(3'd2)))));
  localparam signed [4:0] p16 = ((-2'sd1)<(5'sd12));
  localparam signed [5:0] p17 = (^(&{4{{1{(-3'sd2)}}}}));

  assign y0 = ((p2&&p11)>>>(!a1));
  assign y1 = (-4'sd5);
  assign y2 = ((~&({{2{b1}}}==={(-a4),{a2,b4,a2}}))&(|{(~&(!(-a5))),{(!{p8,p7,p8})}}));
  assign y3 = {($unsigned({$unsigned(b4),(p7<<<b5),(b3&&p1)})>>>{(&{(-{p11,a5,a5})})})};
  assign y4 = $unsigned(((($unsigned(p5)&(p8||p13))>=((b0==p11)>>(b3)))>={1{({1{(p7&p11)}}-(!(p3|p10)))}}));
  assign y5 = (p3<<p16);
  assign y6 = (~&p2);
  assign y7 = (~^(~^(~^(~^{4{(|(~|p3))}}))));
  assign y8 = (((a5&&a5)>>>(b5&b5))!==(-{1{(a2?a2:a3)}}));
  assign y9 = ((~^(((~^{3{b2}})^{3{p3}})))==(-{3{{4{p15}}}}));
  assign y10 = (&(!(~|a5)));
  assign y11 = ((&{1{((a2^~b4)>>{2{a5}})}})>>>((5'd2 * (b0&a2))<<((a1>=b4)<<<(a3>>b0))));
  assign y12 = (!(5'd4));
  assign y13 = ({2{{4{p6}}}}?{3{(~^p4)}}:(~&(~&{(p9?a4:p15)})));
  assign y14 = (5'd17);
  assign y15 = (3'sd1);
  assign y16 = (~|$signed(p3));
  assign y17 = (4'sd1);
endmodule
