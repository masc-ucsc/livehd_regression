module expression_00725(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'sd0)?(-4'sd4):(3'sd1))<<<((2'sd0)!=(-4'sd2)));
  localparam [4:0] p1 = {(~|((3'sd0)<(-4'sd4))),{(2'd0),(4'd15),(4'sd4)},((4'd4)?(-5'sd11):(3'd4))};
  localparam [5:0] p2 = (|((5'd15)-(^(((2'sd1)<<<(4'd8))&((-2'sd1)+(5'd20))))));
  localparam signed [3:0] p3 = ((~|(&{4{(-5'sd8)}}))||(({2{(2'sd0)}}===(~(2'd2)))<<(~|((-4'sd2)===(5'd6)))));
  localparam signed [4:0] p4 = (((2'd1)?(2'sd0):(5'd26))?((5'd19)?(4'sd5):(-3'sd1)):((-4'sd3)?(5'sd0):(4'sd1)));
  localparam signed [5:0] p5 = {2{{2{{1{((2'sd0)?(4'd9):(2'sd0))}}}}}};
  localparam [3:0] p6 = ((-4'sd2)===(3'sd3));
  localparam [4:0] p7 = {1{(5'd2 * ((5'd5)===(3'd3)))}};
  localparam [5:0] p8 = (4'd3);
  localparam signed [3:0] p9 = (|(((2'd2)<<<(4'd10))<<(~(~(-4'sd4)))));
  localparam signed [4:0] p10 = (~^(~^(((!(2'd3))||((2'd3)!==(3'sd3)))>>>(((-5'sd10)===(3'd7))+((3'd3)|(-2'sd0))))));
  localparam signed [5:0] p11 = {3{{(-4'sd3),(4'sd2),(4'sd7)}}};
  localparam [3:0] p12 = (-5'sd4);
  localparam [4:0] p13 = (2'd3);
  localparam [5:0] p14 = ((((3'sd3)^~(-3'sd2))?((3'd0)^(-2'sd1)):((3'd4)<<<(2'sd0)))>>>(((5'd21)?(4'sd7):(-5'sd14))!=((4'd9)>=(-3'sd1))));
  localparam signed [3:0] p15 = {{2{(-5'sd8)}},{(5'd3),(4'd15),(-3'sd0)},((-5'sd8)?(2'd3):(3'd1))};
  localparam signed [4:0] p16 = ((2'sd0)^(-3'sd3));
  localparam signed [5:0] p17 = {(((4'd9)===(3'd5))<<<{(2'd3),(2'd2),(5'd24)})};

  assign y0 = {1{({2{(~&(a0<<b1))}}!==$signed($signed(((!{b1,a5,b1})-(~&$signed(b3))))))}};
  assign y1 = ((-3'sd2));
  assign y2 = {2{(~^(!(~(~^b2))))}};
  assign y3 = {4{((b4?a3:a4)<(b5<<p12))}};
  assign y4 = (2'd2);
  assign y5 = (b4>>>p16);
  assign y6 = {3{({1{p11}}&&{1{p0}})}};
  assign y7 = ((a3&&p13)&(a5^a3));
  assign y8 = (~(((b2===b0)?(p6):$signed(b2))?($signed((p1?p13:p2))^~$signed((p10?b4:a1))):((5'd28)&(4'sd3))));
  assign y9 = (~^(^(p2)));
  assign y10 = (^(~{{(~|p12),{p6},(p2|p7)},$unsigned({(+b0),(5'd18)}),(({4{b4}}))}));
  assign y11 = (+(!{(|$unsigned({(-{p15,b1,p7}),(+{$unsigned(p13),{p0,p10,p2}})}))}));
  assign y12 = (~(~({2{(+(!(p11)))}}>>>$signed(($signed({1{p6}})&(a0<<p7))))));
  assign y13 = ((((b2<<p14)^~(a4&a3))>=((a4%b1)*(a5+p10)))&(((a0<<<b2)!==(a3*b4))&((b3/a2)==(a2&p6))));
  assign y14 = (+(~(((p15?b0:a0)<(|(-p9)))^((a2===b2)>(b5?p3:a3)))));
  assign y15 = $unsigned((((~$unsigned($signed(b3)))?{$unsigned(b2),{a5}}:{a4,b0,b0})));
  assign y16 = (3'sd0);
  assign y17 = {$signed((({a3,p15})?(p1?a0:p4):(p11+p17)))};
endmodule
