module expression_00595(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!{4{(^{2{(4'd7)}})}});
  localparam [4:0] p1 = (^({(-4'sd7),(4'd1),(3'sd1)}?(!((3'd1)==(4'd3))):(^(|(3'sd0)))));
  localparam [5:0] p2 = {1{(4'd4)}};
  localparam signed [3:0] p3 = {{(5'd20),(4'sd3),(5'd7)},{(-4'sd7)},{(-3'sd2)}};
  localparam signed [4:0] p4 = ((|{(^(4'd5)),((-5'sd4)<<(5'd7)),((2'd3)>(-5'sd11))})^({(2'd2),(3'd1)}^{(2'd1),(3'sd3),(-3'sd0)}));
  localparam signed [5:0] p5 = (~(&((~|((2'd3)&(4'd7)))===(+((-4'sd5)-(-3'sd0))))));
  localparam [3:0] p6 = ((3'd4)?{4{(3'd4)}}:(|(2'd0)));
  localparam [4:0] p7 = {(((~|(-3'sd2))===((4'd1)!=(5'd13)))>{(~^(4'd2)),((2'sd0)<(3'sd3))})};
  localparam [5:0] p8 = {4{(5'd26)}};
  localparam signed [3:0] p9 = ((-(&(^{(-4'sd0),(-3'sd2),(5'sd13)})))^(^(5'sd6)));
  localparam signed [4:0] p10 = ((+(5'sd14))>>(3'sd1));
  localparam signed [5:0] p11 = (4'd10);
  localparam [3:0] p12 = {((5'sd14)|(2'sd1)),(5'd23)};
  localparam [4:0] p13 = ({(2'sd1),(-4'sd1),(-3'sd3)}-((2'd2)<<(2'd1)));
  localparam [5:0] p14 = (+(!(-4'sd1)));
  localparam signed [3:0] p15 = ((-(~|(-3'sd3)))?{4{(-2'sd0)}}:(~&(-(4'd0))));
  localparam signed [4:0] p16 = ((~((5'sd15)?(4'sd5):(2'd1)))===(((-4'sd1)^~(2'd3))<<((3'd2)<=(3'd7))));
  localparam signed [5:0] p17 = {1{((3'd6)?(-3'sd3):(2'sd0))}};

  assign y0 = (p2<<<p11);
  assign y1 = (~|p15);
  assign y2 = {(a1?a0:b5),(~|{p2,p0}),{(p10?p10:b0)}};
  assign y3 = {({p1,p17})};
  assign y4 = ((^p14)?(~p7):(-b5));
  assign y5 = (5'd9);
  assign y6 = $unsigned(({(5'd2 * b2),(2'd2),(a4<<a5)}|(~^(!({a5}<(a2<=b5))))));
  assign y7 = ((p9<<a1)<<$signed(p0));
  assign y8 = ($unsigned(($signed((~|b1))>>>$unsigned((~^a1))))==$signed(((^(5'd5))-(^(3'd5)))));
  assign y9 = {4{{p4,p15,p8}}};
  assign y10 = {{({p6}?{p5}:(p0?p5:b4))},{(p9?a1:a5),{p13,p10,p10},{b1,p15,p12}}};
  assign y11 = {b1,b2};
  assign y12 = {(&(-2'sd0)),{p17,p10,p2},(!(-2'sd1))};
  assign y13 = ((a2%a0)%b0);
  assign y14 = ({(b0!==a4),(p4^b2),(a4!=p3)}>>(5'd20));
  assign y15 = (~^(4'sd1));
  assign y16 = (-(+(2'd2)));
  assign y17 = ((a1^~b1)^(a4>=a2));
endmodule
