module expression_00030(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+{{3{((3'sd2)<<<(5'sd8))}},(-2'sd0)});
  localparam [4:0] p1 = {1{(((4'd4)>=(5'd20))?((3'd6)-(5'd17)):((5'd7)&&(3'd5)))}};
  localparam [5:0] p2 = (~&(3'd7));
  localparam signed [3:0] p3 = {1{{(-3'sd0),(5'd30),(3'd6)}}};
  localparam signed [4:0] p4 = {2{{{1{((4'd10)<(4'sd3))}},((2'd3)|(3'd1))}}};
  localparam signed [5:0] p5 = (((3'sd1)&&(3'd7))>((5'd18)>=(3'sd0)));
  localparam [3:0] p6 = {(~(&{(5'd2 * {((5'd23)^(2'd1))})}))};
  localparam [4:0] p7 = ((-4'sd2)?(+(2'sd0)):(2'd2));
  localparam [5:0] p8 = {{1{((4'sd3)?{3{(2'd2)}}:{3{(2'd1)}})}},{4{{(3'd5)}}}};
  localparam signed [3:0] p9 = ((-3'sd0)?(2'd0):(-2'sd0));
  localparam signed [4:0] p10 = (^((~(~|(&(|(-5'sd8)))))<((-5'sd4)===(~(-5'sd5)))));
  localparam signed [5:0] p11 = (3'd6);
  localparam [3:0] p12 = {2{{(~(2'd3)),(&(2'sd0)),{(-2'sd1),(4'd10),(-3'sd0)}}}};
  localparam [4:0] p13 = (((5'd2)<(2'd1))&&{(2'sd0),(5'd28)});
  localparam [5:0] p14 = ((-3'sd2)/(4'd4));
  localparam signed [3:0] p15 = (((!(2'sd0))!==(~(3'd5)))>((~^(3'sd3))!=((4'd7)-(2'd0))));
  localparam signed [4:0] p16 = (|(((5'sd7)<(3'd5))>((-4'sd5)|(-3'sd0))));
  localparam signed [5:0] p17 = (2'd3);

  assign y0 = ((~((&(a3/b1))/a0))&&(+(-(&(b2>p17)))));
  assign y1 = (($unsigned((-4'sd3))>>>(b1|a4))===$signed($unsigned(((b4&b2)<<<(2'sd1)))));
  assign y2 = ((a0===b3)||(a0?a5:a4));
  assign y3 = (^(~^(~&(~&(^(4'd5))))));
  assign y4 = (~|$signed(((p1?p12:p1)?{b3,b0,p17}:({p3}<(~^p16)))));
  assign y5 = (2'd1);
  assign y6 = ((((b0!=a5)^~{b0,b0,b2})&&((a3>b3)&(a3>>>b4)))+{(((a0===b4)!==(a4|a5))-({b1}|{b1,a4}))});
  assign y7 = (~^($signed(p0)?{p3,p11}:$signed(b1)));
  assign y8 = (a0||a2);
  assign y9 = ({1{p9}}?(p15==b3):(a0!==a2));
  assign y10 = (p8?b2:b5);
  assign y11 = (-3'sd2);
  assign y12 = (~^(-(+(({p9,p15}>>>(p0^~p11))+(|(-{p4,b2}))))));
  assign y13 = (-4'sd7);
  assign y14 = {(~^a4),(+b3)};
  assign y15 = (((-3'sd1)-(2'd3))?((b0!==a2)?(3'd6):(-3'sd2)):(2'd3));
  assign y16 = (~(-4'sd4));
  assign y17 = (p8?a2:a0);
endmodule
