module expression_00147(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~|(((5'sd11)+(-5'sd1))%(-2'sd1)))<=(^(((2'd2)>(5'd21))||((3'd5)%(2'd2)))));
  localparam [4:0] p1 = {3{{1{{4{(5'd14)}}}}}};
  localparam [5:0] p2 = (~|(-(!(+(~(^{{{{4{(~(-3'sd2))}}}}}))))));
  localparam signed [3:0] p3 = (~{{(~^(!((-3'sd0)>>>(-5'sd6))))},{(~|(3'd4)),{1{(-5'sd14)}},(&(5'sd2))}});
  localparam signed [4:0] p4 = (&((((3'd3)>>(-3'sd2))?((2'd2)<<(-2'sd0)):((5'd1)/(3'd6)))<<((^(|(2'd3)))/(5'sd7))));
  localparam signed [5:0] p5 = (((((4'sd6)>=(2'd1))<<((5'sd7)<<<(5'd2)))^(6'd2 * ((2'd0)<(4'd6))))>=((((-3'sd3)>=(2'd3))!==((3'sd0)&&(3'd0)))>=(4'd2 * (6'd2 * (3'd1)))));
  localparam [3:0] p6 = (({(5'd7),(2'd3),(4'd0)}||{4{(2'd3)}})!==((3'sd1)=={(3'd1),(4'd7)}));
  localparam [4:0] p7 = (^(-4'sd2));
  localparam [5:0] p8 = ((!(3'd1))!==(+(4'd8)));
  localparam signed [3:0] p9 = ({3{(5'sd1)}}+(((5'd30)<=(4'd8))<((5'sd0)^~(-5'sd13))));
  localparam signed [4:0] p10 = {(3'd2),(-3'sd1),(5'sd7)};
  localparam signed [5:0] p11 = (-{{{(-5'sd5)},{(4'd15),(5'sd12)},(~|(3'd4))},{(5'd2 * (5'd1)),{(-3'sd3),(3'sd1)},(!(-4'sd7))}});
  localparam [3:0] p12 = (6'd2 * ((3'd7)|(4'd13)));
  localparam [4:0] p13 = ((~^(&(5'd16)))==({2{(3'sd3)}}|(~|(-5'sd3))));
  localparam [5:0] p14 = {2{(5'd24)}};
  localparam signed [3:0] p15 = (((~^{3{(-2'sd0)}})>>>(!{(2'd0),(4'd15)}))>>>{4{(-(4'd15))}});
  localparam signed [4:0] p16 = ((((-5'sd11)&&(5'd24))!==(|{(-4'sd2),(3'd0)}))<=((~|(+(4'd10)))>((5'd20)?(3'sd1):(5'd8))));
  localparam signed [5:0] p17 = (~^(((5'd18)^~(5'd0))^~(!((-2'sd0)?(5'd3):(5'd28)))));

  assign y0 = (|((((p4||p4)<<<(p0^p7))!=(!(p1<<p11)))>>(((p10>>>p2)<=(p17-a4))^~(-(p11>>p7)))));
  assign y1 = $signed((((p5&p10)?(p13?a0:b5):(-3'sd0))?({b0,p16,b3}>={b2}):{{p17,p13,b3},(6'd2 * p14)}));
  assign y2 = (~|(p9?p16:p11));
  assign y3 = ((~|(~^(2'sd1)))?{3{(2'd1)}}:{1{(4'd6)}});
  assign y4 = (4'd15);
  assign y5 = {2{(p3?p16:p17)}};
  assign y6 = {{4{p0}}};
  assign y7 = (5'sd0);
  assign y8 = (a0?p7:p14);
  assign y9 = (((a0?b5:a2)-(a2?b3:a5))?((p4>>>p2)>=(a1?b2:a0)):((b3?b4:b0)?(p3^p17):(b2?a4:b4)));
  assign y10 = (-5'sd10);
  assign y11 = ({{4{b0}},{2{b2}},{p2,p13,p0}}?({3{b3}}?(b1?b1:a3):{p8,a0}):{{4{a3}},(~&p5),(p14?p14:b4)});
  assign y12 = ((-5'sd15)^(5'sd14));
  assign y13 = {2{({(p14-p9)}|(&{2{p11}}))}};
  assign y14 = {((~&p15)|(~a3))};
  assign y15 = ({((a0?a5:b2)>>(a2==a1))}<{$unsigned($unsigned((b1?a0:b2)))});
  assign y16 = ((((b2?a3:b1)?(a1>>>a1):(~a2))^((b3?b5:b2)?(!b2):(b5?b0:b1)))===(+(&(&((&b4)?{1{b1}}:(b4>>a3))))));
  assign y17 = (+(b5^~b1));
endmodule
