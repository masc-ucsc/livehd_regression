module expression_00790(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(3'd7));
  localparam [4:0] p1 = {(3'd3),(3'd5),(2'd0)};
  localparam [5:0] p2 = ((~&(((4'sd3)<=(3'sd1))+{2{(4'd4)}}))-(((2'sd1)&&(4'd0))===((2'd3)<(4'd9))));
  localparam signed [3:0] p3 = ({((-5'sd12)?(4'sd4):(3'sd3))}?{(3'sd2),(5'd26),(3'sd3)}:((5'sd6)?(2'd3):(4'sd4)));
  localparam signed [4:0] p4 = ((&(3'd5))?((5'd2)?(4'd5):(-5'sd5)):((3'd5)?(2'd0):(-5'sd12)));
  localparam signed [5:0] p5 = (((-4'sd5)?(3'd6):(5'sd12))?{(4'sd6),(5'sd6),(4'sd1)}:((-5'sd1)<=(3'sd1)));
  localparam [3:0] p6 = {{4{(3'sd1)}},(~^(2'd0)),((5'd12)&&(-2'sd1))};
  localparam [4:0] p7 = (((5'd16)<(5'd25))/(-4'sd4));
  localparam [5:0] p8 = (-4'sd6);
  localparam signed [3:0] p9 = {{(2'd3)},{(4'd4)},(6'd2 * (3'd7))};
  localparam signed [4:0] p10 = (((-3'sd1)/(-3'sd1))*(-((5'sd5)*(3'd6))));
  localparam signed [5:0] p11 = ({((3'd6)<=(3'd7)),(4'd5),{2{(4'd7)}}}<<<{((3'd0)^(3'sd3)),{(2'd3)}});
  localparam [3:0] p12 = (&(-4'sd7));
  localparam [4:0] p13 = {2{{(+{2{(2'sd0)}})}}};
  localparam [5:0] p14 = ({3{(-3'sd3)}}<<<({2{(-5'sd8)}}!==(2'd1)));
  localparam signed [3:0] p15 = {1{(!{4{(((-5'sd9)|(-4'sd7))^(~^(4'sd2)))}})}};
  localparam signed [4:0] p16 = (~|(+(!(~&(-(~|(-(+(^(+(^(!(!(~(5'd4)))))))))))))));
  localparam signed [5:0] p17 = ({{(-4'sd1)},{(4'd4),(3'd3)},{(3'sd1)}}>>(((5'd29)&(-3'sd2))>=((3'd2)^(4'd12))));

  assign y0 = {(({b4,a0,a1}==={(a0==b4)})|((a4>>>a1)>={(a4^a1)}))};
  assign y1 = {3{{1{(^{4{p17}})}}}};
  assign y2 = (p0?p4:p5);
  assign y3 = ((p5?p3:a1)?(a4==p10):(b1!==a0));
  assign y4 = (((^b3)?(~&a3):(-a0)));
  assign y5 = (+(4'd2 * (a1!==b1)));
  assign y6 = (a1?a0:a2);
  assign y7 = (-{(|(-((^((|(-b1))|(-{3{b5}})))!=={3{(+a4)}})))});
  assign y8 = {(!(^(p12?a2:p10))),(b5?b0:p8),(&(^(^p1)))};
  assign y9 = {4{{a0,a0,b5}}};
  assign y10 = $signed({(~|(&(a5|b5)))});
  assign y11 = ({{({3{{p13,p11}}})}}&&($signed(((p14<p9)>$unsigned(p10)))<<<{{p5,p16,p10},{p5,a4},(p15-p6)}));
  assign y12 = ({1{{1{((&(a2?a1:p2))?{a4,p12}:(p1?p10:p6))}}}}|((b4===a0)?(~{p10}):(a0==p16)));
  assign y13 = (-2'sd0);
  assign y14 = (4'd2 * (5'd26));
  assign y15 = ({2{(5'd2 * (&(p2<<<p0)))}}>>((~&({3{p3}}|(b3-b2)))>=((b2===a1)^(p5||p1))));
  assign y16 = (-3'sd1);
  assign y17 = {{b3,p12,a5},((b5?p2:p4)^(b1-p2)),(5'd28)};
endmodule
