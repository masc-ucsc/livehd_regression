module expression_00248(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'sd1);
  localparam [4:0] p1 = (((5'd12)>>(2'd2))?{3{(2'sd0)}}:(4'd7));
  localparam [5:0] p2 = (((!(4'sd0))?((2'd3)>=(2'sd0)):(3'd1))!==(-4'sd3));
  localparam signed [3:0] p3 = ((2'sd0)!=(3'd4));
  localparam signed [4:0] p4 = ({(4'd3),(-5'sd12)}?((3'd5)?(-3'sd3):(4'sd5)):(~&(~|(5'sd12))));
  localparam signed [5:0] p5 = (^(~|(-(!(+(&(~|(|(~^(|(!(~&(3'd5)))))))))))));
  localparam [3:0] p6 = (3'sd3);
  localparam [4:0] p7 = (6'd2 * (~(4'd2)));
  localparam [5:0] p8 = (-5'sd13);
  localparam signed [3:0] p9 = (4'd14);
  localparam signed [4:0] p10 = (2'd1);
  localparam signed [5:0] p11 = (((4'd1)?(2'd3):(-5'sd3))?{2{(3'd6)}}:{1{(3'd3)}});
  localparam [3:0] p12 = ({((2'd3)?(2'd1):(4'sd7)),(!(5'sd14)),(~&(4'd1))}||(6'd2 * ((2'd0)?(4'd15):(5'd25))));
  localparam [4:0] p13 = ((5'd2 * (2'd3))?(3'd4):((2'sd1)?(4'd6):(3'sd3)));
  localparam [5:0] p14 = (^(((-4'sd3)<<(2'd1))!==(-2'sd0)));
  localparam signed [3:0] p15 = (2'd1);
  localparam signed [4:0] p16 = (3'sd1);
  localparam signed [5:0] p17 = {4{{(4'sd4),(5'd8),(-5'sd10)}}};

  assign y0 = $unsigned((5'd15));
  assign y1 = ($signed((a3?b1:p16))?(a1||a3):(~(p17|a0)));
  assign y2 = $signed((+(($unsigned((!$signed(($unsigned(((p12<<<p6)<(a2>>>p1)))==(&$unsigned((~|(p8))))))))))));
  assign y3 = {3{(a2?p17:p11)}};
  assign y4 = (~|(~&(-{1{(~&((b3||b3)+(~&b4)))}})));
  assign y5 = ((+a1)<<(~b1));
  assign y6 = {1{({1{(^{4{b2}})}}===((~^a1)>={1{b1}}))}};
  assign y7 = {4{p2}};
  assign y8 = ({((p7<p10)),{4{p16}},{p2,p8,p13}});
  assign y9 = {((&a3)||(+p2)),((-2'sd0)&(b5+a2)),(&(-4'sd1))};
  assign y10 = {$signed((a2>>>b3))};
  assign y11 = ((b0?a3:a3)?(-2'sd1):(b0?a3:b5));
  assign y12 = (-(b4));
  assign y13 = (~&{(5'd2 * p6),(p8&p7),(p9&p17)});
  assign y14 = ((~|(~(b2?b4:p10)))?(~(&(&(p13==b2)))):((|b5)^~(a4?a2:p6)));
  assign y15 = (-5'sd1);
  assign y16 = (((|{b0,a4})?$unsigned((b4<=p5)):(&(!(|b0)))));
  assign y17 = (5'd2 * {1{(p6!=a1)}});
endmodule
