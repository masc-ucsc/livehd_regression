module expression_00830(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(2'd0));
  localparam [4:0] p1 = (4'd2 * ((2'd3)<<(2'd1)));
  localparam [5:0] p2 = {2{{(&{1{(4'sd5)}}),{4{(5'd19)}}}}};
  localparam signed [3:0] p3 = (~(&(~&(!(((3'd3)==(-2'sd1))&&(|(5'd23)))))));
  localparam signed [4:0] p4 = (((~&((-5'sd5)!=(5'd18)))+(((5'd31)^(5'sd6))<(~(-5'sd0))))>=(4'sd2));
  localparam signed [5:0] p5 = {1{(4'sd5)}};
  localparam [3:0] p6 = (((-4'sd1)?(-2'sd1):(2'd2))^~(3'd3));
  localparam [4:0] p7 = ({((4'sd1)!==(4'd14)),((5'd17)?(-3'sd0):(5'd26))}|{(3'd1),(2'd1),(4'd8)});
  localparam [5:0] p8 = (~|(~|(-2'sd0)));
  localparam signed [3:0] p9 = ((!((^{(3'd6)})||{(2'd3),(4'd14)}))==(&{(((-5'sd1)-(-4'sd3))?(^(4'd6)):{(-2'sd1),(4'd4),(5'sd3)})}));
  localparam signed [4:0] p10 = ((4'd13)<<(-3'sd0));
  localparam signed [5:0] p11 = ((-2'sd0)?(3'sd3):{4{(3'sd0)}});
  localparam [3:0] p12 = ((3'd7)?(5'd1):(5'd13));
  localparam [4:0] p13 = {(~{({(3'd1),(-3'sd3)}>=(-5'sd3))}),{((5'd18)>=(2'd3)),(^{(3'sd0)})}};
  localparam [5:0] p14 = (+(((-4'sd5)?(5'sd10):(4'd13))?{2{(5'd13)}}:((-4'sd3)?(5'sd1):(2'sd1))));
  localparam signed [3:0] p15 = (+(&(+({1{{(5'd18),(3'd7),(-4'sd7)}}}>((&(2'sd0))>>>(+(2'd3)))))));
  localparam signed [4:0] p16 = (~^(~{4{(4'd5)}}));
  localparam signed [5:0] p17 = ((5'sd1)>>(2'd0));

  assign y0 = {(!{({1{(~{p4})}}>>(p3?p15:p10))})};
  assign y1 = (2'sd0);
  assign y2 = (&(-{4{(5'd2 * {3{p2}})}}));
  assign y3 = ($unsigned(((b3?a3:p4)?{b0}:(b0?a4:b2)))?((5'd2 * p6)?(a4?a3:a0):$unsigned(a1)):{(b0<<<a3),(a2?a1:p2)});
  assign y4 = (+(-{{{b4,a5,b4},(+{b3,b5,a1})},{(~((^(~&b5))&(a3&a2)))}}));
  assign y5 = $signed((a1>p16));
  assign y6 = (~&(-(!(((p11?b1:p17)?(p10?p5:a2):{2{p6}})>>>((~^a5)?(|a5):(a1!=a4))))));
  assign y7 = ({{((p3>>p0)>={4{a3}}),(5'd2 * (!p14))}}&(((b5>>a4)-(!b4))==={4{b0}}));
  assign y8 = {{4{p9}}};
  assign y9 = {2{{3{{a1}}}}};
  assign y10 = (b2?p6:p0);
  assign y11 = (!(|(~(({a4,a3}!==(b4<=b4))>>({b4}<<(a0^~a5))))));
  assign y12 = ((((a3+a0)>>>(^a1))||($signed(b0)<<<{3{a3}}))=={{(a5?b3:b4),((b3|b2)),{a3,a2,b0}}});
  assign y13 = (((p2>p13)*(a1===b1))^((p5*p4)>>>(p12>>p12)));
  assign y14 = $unsigned((|({p3,a0}?(p17+a1):$unsigned((~&p9)))));
  assign y15 = {2{(a1>>b4)}};
  assign y16 = ({2{p2}}?{3{p11}}:(p9&&p17));
  assign y17 = ($signed(((2'd1)<<(5'd6)))||($signed($signed(b4))!=(p6||b5)));
endmodule
