module expression_00231(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(~(~^(&((4'd15)|(2'd2))))));
  localparam [4:0] p1 = {{{(5'd12),(2'sd0)}},{{(2'd1),(3'd0),(2'd2)},{(-5'sd3),(3'sd2)}},((~|(3'd3))+{(3'd5)})};
  localparam [5:0] p2 = {((|(3'd3))!==(-(-3'sd3)))};
  localparam signed [3:0] p3 = (({((5'd4)!==(5'd27))}==(~{3{(3'sd1)}}))|{(6'd2 * (5'd16)),((-2'sd1)!==(3'd2))});
  localparam signed [4:0] p4 = {(5'd5),(-4'sd7),(-4'sd1)};
  localparam signed [5:0] p5 = (4'sd2);
  localparam [3:0] p6 = (({3{(-5'sd13)}}<((2'd1)<<(-5'sd5)))?(((3'd5)-(4'd5))?{1{(2'd3)}}:{1{(-2'sd0)}}):(((3'd2)&&(3'd5))&&((3'sd1)<=(-3'sd0))));
  localparam [4:0] p7 = ((-2'sd0)/(3'd7));
  localparam [5:0] p8 = {4{(-2'sd1)}};
  localparam signed [3:0] p9 = (3'd5);
  localparam signed [4:0] p10 = (^(!((3'd1)!==(-2'sd1))));
  localparam signed [5:0] p11 = ({1{{1{{4{(5'sd1)}}}}}}|(((3'd2)<(4'd7))?((3'd6)===(2'sd0)):{3{(2'd3)}}));
  localparam [3:0] p12 = ((((3'sd0)?(2'sd1):(4'sd6))!=={(5'd15),(3'd6),(-2'sd0)})^~{((-3'sd0)>(2'd0)),((5'sd0)?(5'sd2):(-3'sd1)),((4'd11)?(2'd0):(2'd2))});
  localparam [4:0] p13 = (5'sd14);
  localparam [5:0] p14 = ((&{{(&{(-5'sd2),(-4'sd6),(3'd2)})}})==({(3'd7),(4'd11)}<<<((3'd5)-(5'd15))));
  localparam signed [3:0] p15 = ((-2'sd0)==(4'sd6));
  localparam signed [4:0] p16 = ((~&((-5'sd7)<(5'd4)))||((-5'sd0)?(2'sd1):(-5'sd1)));
  localparam signed [5:0] p17 = (!(^((~&((3'd7)%(-3'sd0)))/(2'd0))));

  assign y0 = (a3?b2:a0);
  assign y1 = (2'd2);
  assign y2 = (5'd25);
  assign y3 = (|$unsigned((p13?a4:p14)));
  assign y4 = ((!(-$signed(((~&p9)^~$signed(p12)))))>>($unsigned($signed((p14)))==$unsigned((p14<p4))));
  assign y5 = (&(((3'd1)>>(b0!==b1))-(5'd10)));
  assign y6 = (~|{2{{{3{a3}},{p11,a2,b2}}}});
  assign y7 = {{4{{b2,b5,b2}}},((b0^~b4)<=$signed({3{a3}}))};
  assign y8 = $unsigned((((~|(+(3'sd2)))||((-4'sd5)>>$unsigned(b5)))));
  assign y9 = (~&(-((^((~^p0)&&(&p16)))+((~|b0)>(a5>=b4)))));
  assign y10 = (-(((^(a3?p11:p10)))<<((p13>>b2)?(3'd1):(p12?p7:a2))));
  assign y11 = (((((b4^~b0)^~$signed(b1))>((a2/b0)%a2)))==$signed((((b1<<b0)&(b3!==b2)))));
  assign y12 = ((3'sd2)?{b2,a5,b2}:(5'd2 * {p7,b0,a0}));
  assign y13 = (~(+((b3?p16:p13)?{4{p0}}:(|a1))));
  assign y14 = (({a1}?(b2):(a5?a5:a1)));
  assign y15 = (^(~|(~(~^p6))));
  assign y16 = (-{({b1,b5,p3}-((p1?p6:b2)|(|p10))),((+(b2&p6))>=(b2?p10:b0))});
  assign y17 = (((p14?p6:a1)!=(^p2))-((p8>p6)>=(p12||p13)));
endmodule
