module expression_00249(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({2{{3{(-4'sd2)}}}}+(((3'd3)&(5'd18))?((-4'sd3)>(-4'sd6)):{2{(2'sd1)}}));
  localparam [4:0] p1 = {4{{1{((2'd3)<<(4'd13))}}}};
  localparam [5:0] p2 = ((~&(5'sd15))?(|(4'd11)):(~&(-4'sd6)));
  localparam signed [3:0] p3 = (~|(|(5'd6)));
  localparam signed [4:0] p4 = (-3'sd1);
  localparam signed [5:0] p5 = ((5'd25)?(~&(4'd7)):(-(-2'sd0)));
  localparam [3:0] p6 = {{((3'd1)?(-3'sd1):(2'd2)),(|(5'd2))}};
  localparam [4:0] p7 = (5'd9);
  localparam [5:0] p8 = (-((~(~&{2{((2'd3)^~(-2'sd1))}}))<<(((-2'sd1)|(-5'sd15))&&{3{(3'd2)}})));
  localparam signed [3:0] p9 = (({2{(3'd0)}}^((4'd13)==(4'd8)))?(+(-((-3'sd2)>(-4'sd4)))):((|(3'd2))<<<{(-2'sd1),(4'd6),(-4'sd6)}));
  localparam signed [4:0] p10 = {(2'd1),{((2'd2)|(3'd6)),(~|(-3'sd0))}};
  localparam signed [5:0] p11 = (((5'd3)|(2'd0))?(-4'sd5):((3'd1)>(5'd31)));
  localparam [3:0] p12 = ((|(^(3'd0)))?((5'd0)?(-4'sd4):(-3'sd2)):((5'd22)||(5'd4)));
  localparam [4:0] p13 = (3'sd1);
  localparam [5:0] p14 = ({{(3'sd2),(3'd7)}}?(((3'd0)<<(-4'sd0))<=((-5'sd6)?(2'd2):(3'sd3))):(~|{3{(3'd7)}}));
  localparam signed [3:0] p15 = {(&({(2'd0),(3'sd1),(4'sd7)}&&(+((4'd7)?(-3'sd2):(5'd5))))),((~{(2'd2),(-4'sd1)})?(+(~(2'd3))):(^((4'd5)<=(3'sd0))))};
  localparam signed [4:0] p16 = ((4'd1)+(^((2'd2)&(-5'sd11))));
  localparam signed [5:0] p17 = (5'd2 * {(5'd20),(2'd3),(4'd12)});

  assign y0 = (p1?b2:p14);
  assign y1 = {4{{2{{3{a5}}}}}};
  assign y2 = (^(+{{(~^(p5^~p16))},{p17,a0,p2}}));
  assign y3 = (p0?a1:a5);
  assign y4 = (((a1>a4)!=={3{a2}})-((-2'sd1)!=(a4<=a0)));
  assign y5 = (({4{a2}}&&(~&(a3?b5:a0)))^~(^{{4{a3}}}));
  assign y6 = (b5?b1:p12);
  assign y7 = (-2'sd0);
  assign y8 = {({((p6?p5:b2)==(2'd1)),(({p10,p12}+($signed(b3))))})};
  assign y9 = (!(~{4{{1{(&a0)}}}}));
  assign y10 = (((a4/b3)==(a0|p11))<=((b2&&b1)|(~^(-5'sd7))));
  assign y11 = {1{b3}};
  assign y12 = (((p2&b1)/p3)?((p16<<<p9)?(p5>>p3):(p5!=p9)):((b3?a2:p2)?(p13<<p15):(p0||b1)));
  assign y13 = (p3!=p4);
  assign y14 = (2'sd0);
  assign y15 = $unsigned((-2'sd0));
  assign y16 = ({3{(5'sd12)}}+((p12<=p3)>(~^(p13>p15))));
  assign y17 = (p12<<<p6);
endmodule
