module expression_00441(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(5'd16),((-2'sd1)?(-3'sd2):(3'sd0))};
  localparam [4:0] p1 = (((-5'sd13)?(3'sd3):(4'sd1))||(2'd1));
  localparam [5:0] p2 = ((3'd0)!==(((-5'sd6)?(4'd4):(4'd11))!=((3'd7)&(3'd2))));
  localparam signed [3:0] p3 = (2'd0);
  localparam signed [4:0] p4 = ((3'sd0)>(-4'sd5));
  localparam signed [5:0] p5 = {(2'd2),(5'sd1),(2'd2)};
  localparam [3:0] p6 = {(((5'd12)==(5'd23))^~(!(-3'sd0)))};
  localparam [4:0] p7 = {(4'd11)};
  localparam [5:0] p8 = {4{(2'd3)}};
  localparam signed [3:0] p9 = {4{({2{(-3'sd0)}}<((-5'sd6)<=(4'd4)))}};
  localparam signed [4:0] p10 = ((2'sd0)>(3'sd0));
  localparam signed [5:0] p11 = {({2{(2'd0)}}?((3'd6)?(3'sd3):(4'sd2)):((-4'sd5)?(2'd3):(-5'sd15)))};
  localparam [3:0] p12 = ({(3'd0),(5'sd15),(5'd24)}^~{3{(5'd10)}});
  localparam [4:0] p13 = ({(2'd3)}>>>(4'd0));
  localparam [5:0] p14 = (4'd2);
  localparam signed [3:0] p15 = (2'sd0);
  localparam signed [4:0] p16 = ((-4'sd0)^~((-4'sd7)<=(-3'sd2)));
  localparam signed [5:0] p17 = {(+(~|((3'd6)<=(2'sd1)))),(((4'sd2)<=(3'd0))<((3'sd1)?(-2'sd0):(-5'sd0))),{((2'sd0)||(4'sd1)),((5'd8)|(-2'sd0))}};

  assign y0 = (((~(-4'sd3))||{4{a5}})+((~|(+b1))+(b2^p10)));
  assign y1 = (4'sd2);
  assign y2 = {{{{4{b0}}}},(5'd30),{(2'd1),(b3^~b3)}};
  assign y3 = ((&(-(5'sd6)))^~(!$signed((4'd1))));
  assign y4 = (2'sd0);
  assign y5 = (((b0==b5)>={3{a5}})===(5'd2 * (4'd12)));
  assign y6 = (((p12<<<a0)?(3'd0):(+a4))^(4'd13));
  assign y7 = ((p5|b2)>(a4&a0));
  assign y8 = ({$signed({p17,p7,p6}),{p16,p11,p12}}>(~((!(p15>=a5))<<({p3,p7}<=(a3===b1)))));
  assign y9 = {1{$unsigned((3'sd2))}};
  assign y10 = ((~|(a0?b5:a5))?(b3?b5:a2):((b5||a2)^(~&a0)));
  assign y11 = ((b2?b3:p11)>={2{p13}});
  assign y12 = ({{p11,p16,p4},{2{p2}}}<<<(+{3{{3{p1}}}}));
  assign y13 = (($signed((p13%a3))-(a2-a1))>>(-3'sd3));
  assign y14 = (3'd4);
  assign y15 = (-3'sd2);
  assign y16 = ((b5>>>p15));
  assign y17 = {1{((!(&b5))?(-3'sd1):{2{b3}})}};
endmodule
