module expression_00386(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd0);
  localparam [4:0] p1 = (~^{({(3'sd1)}<(~(4'sd3))),{(!(-5'sd11)),((5'sd7)<<(2'sd1))},(((4'd4)<(2'd2))!={(3'd5),(-3'sd0),(4'sd0)})});
  localparam [5:0] p2 = (((-5'sd7)?(3'd5):(4'd5))?((4'd3)+(-5'sd11)):((3'd2)?(3'd1):(-3'sd1)));
  localparam signed [3:0] p3 = (+(((4'sd0)?(-4'sd2):(4'd13))?{(2'd3),(5'd15),(5'sd5)}:(~^(-4'sd5))));
  localparam signed [4:0] p4 = (5'd1);
  localparam signed [5:0] p5 = ({4{(5'd14)}}==({(4'd13),(-4'sd5)}!={2{(3'd4)}}));
  localparam [3:0] p6 = (({2{((2'sd0)?(3'd2):(5'd16))}}<<((2'sd1)?(-3'sd0):(-3'sd1)))^~{1{((~&(-2'sd1))?((-5'sd10)-(4'd6)):(~&(3'd7)))}});
  localparam [4:0] p7 = ({1{(-4'sd6)}}<((2'sd0)>=(2'd2)));
  localparam [5:0] p8 = ((((2'sd0)-(2'sd1))?(^(2'sd1)):(-(-5'sd4)))||((~&(5'sd14))>>(&(-5'sd10))));
  localparam signed [3:0] p9 = ((-(2'sd1))?(+(3'd4)):((3'sd0)?(-3'sd2):(4'd4)));
  localparam signed [4:0] p10 = (6'd2 * {3{(5'd6)}});
  localparam signed [5:0] p11 = {1{({3{(+(3'sd0))}}==={{(3'd7),(-5'sd11),(4'sd4)},((3'sd0)^~(3'sd1)),{1{(4'sd2)}}})}};
  localparam [3:0] p12 = ((3'sd3)>>(-3'sd1));
  localparam [4:0] p13 = (((4'd4)-(-3'sd3))^~{3{(3'd6)}});
  localparam [5:0] p14 = {4{(5'd27)}};
  localparam signed [3:0] p15 = {3{(4'd3)}};
  localparam signed [4:0] p16 = (-3'sd2);
  localparam signed [5:0] p17 = {{3{((3'sd1)||(-5'sd11))}},(-(((4'd8)<<(4'd11))<{4{(4'd10)}}))};

  assign y0 = (($unsigned(p2)<<<(p2+p8)));
  assign y1 = {4{{3{p7}}}};
  assign y2 = (((p1?p15:a0)?(p14?a5:b0):(p5?p11:p15))?((p11*a0)?(!p13):(4'd13)):((p6<=p2)>=(-3'sd1)));
  assign y3 = (~&(3'd3));
  assign y4 = ($signed(({4{b0}}&(p7?b2:a4)))^~(-((p6>>p2)&&(b1?a5:a2))));
  assign y5 = ($signed(({p10,b4,b0}<<<(b3!==b3)))!=(-({(b1)}^(a3?p16:b0))));
  assign y6 = (4'd6);
  assign y7 = ((((b2<<<a1)!=(a4==b1))||((b4-a2)<(a4<<a4)))===(((a3<=a1)<=(a2^~a2))&((a3==b1)<<<(a3^~b2))));
  assign y8 = {2{{4{a5}}}};
  assign y9 = ({1{{(b5),(6'd2 * b0),{1{a3}}}}});
  assign y10 = ({p1,a0,b2}<=((b4<a0)));
  assign y11 = {(~|{2{{(p0?a3:p14)}}}),(~|(^{(~^(p13?a5:b5))})),{2{{b2,b3,b0}}}};
  assign y12 = (((b0-a5)>>(2'd1))&&({(3'd7)}<<(b3^~b4)));
  assign y13 = (5'sd12);
  assign y14 = (!((!$signed($unsigned($unsigned((^{2{(+a2)}})))))<<{1{{3{{4{p9}}}}}}));
  assign y15 = (((p10?p6:a2)>({b5}>>(p8||p8)))<<{{{p11}},(p0?a4:p12),(a4>>>p3)});
  assign y16 = {1{{4{(4'd7)}}}};
  assign y17 = (~|((|(-{4{b4}}))==={1{(b3?a2:b3)}}));
endmodule
