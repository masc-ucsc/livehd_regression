module expression_00254(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd30)<<(2'sd1));
  localparam [4:0] p1 = ((~|((3'd3)>>>(5'sd5)))&&((3'sd0)?(5'd0):(-2'sd0)));
  localparam [5:0] p2 = (!(~&(2'd0)));
  localparam signed [3:0] p3 = (~|(~(^{((!(!(3'sd3)))>>{(5'd13),(5'sd11),(3'd0)})})));
  localparam signed [4:0] p4 = (~{((2'd2)==(4'd6))});
  localparam signed [5:0] p5 = ({2{(4'sd4)}}?((3'd0)?(4'sd7):(2'd1)):((5'd21)?(-3'sd1):(5'sd6)));
  localparam [3:0] p6 = (|(~(|(~|(!(|{2{(!(~|(3'sd3)))}}))))));
  localparam [4:0] p7 = ((((-3'sd1)<(2'd1))>(~(4'sd3)))?(((2'd3)?(-3'sd1):(4'd9))==(5'd2 * (2'd2))):{4{(2'd2)}});
  localparam [5:0] p8 = (((3'sd2)||(5'd29))<<<((4'd6)||(4'sd6)));
  localparam signed [3:0] p9 = ((|(5'd10))?((2'd1)?(5'd20):(-5'sd2)):((3'd0)>=(-4'sd1)));
  localparam signed [4:0] p10 = {1{(+((^(2'd2))?(^(5'd27)):{4{(4'sd7)}}))}};
  localparam signed [5:0] p11 = (+((|(-4'sd2))?(5'd2 * (4'd4)):((5'sd13)<(2'sd0))));
  localparam [3:0] p12 = {(((3'd3)<<(-4'sd4))+((2'd0)<<<(2'd0))),({(-5'sd14),(-4'sd6),(-2'sd0)}^((3'sd0)^(2'sd0))),({(3'd4),(4'd8),(5'sd0)}||{(4'd5),(3'd1)})};
  localparam [4:0] p13 = ((((-3'sd2)^(-4'sd4))>>(^((5'd18)&(-3'sd2))))>>>{{1{{1{{((-5'sd15)+(4'd14)),{2{(2'd0)}}}}}}}});
  localparam [5:0] p14 = ({(5'sd5)}!={(3'sd1),(5'sd13)});
  localparam signed [3:0] p15 = ((2'd0)===(3'd7));
  localparam signed [4:0] p16 = (((5'sd0)?(-4'sd4):(2'd1))>>((3'sd1)==(3'd5)));
  localparam signed [5:0] p17 = (~&((((-2'sd1)?(3'sd1):(3'sd3))?((3'd3)?(2'd2):(3'd7)):(&(3'sd0)))>>(&(+((3'sd2)||(-4'sd0))))));

  assign y0 = ((b5&a3)%a2);
  assign y1 = (+a3);
  assign y2 = (~{({(2'd1),(|p15)}^(4'd4)),({2{(-5'sd4)}}&&{4{p3}})});
  assign y3 = {2{(^((~b3)?$unsigned(b1):(|b1)))}};
  assign y4 = (+(5'sd2));
  assign y5 = (-4'sd3);
  assign y6 = ((~&(2'sd1))+(2'sd1));
  assign y7 = {2{(((b2&a5)?$unsigned(p11):$unsigned(a2)))}};
  assign y8 = ((b5<<<b3)|(a1^~b2));
  assign y9 = (((p3>>>p12)>={p2,p2,p17})?{{(p6?p13:p8)}}:{(p3?p15:p8),(p0^p7)});
  assign y10 = (6'd2 * (a1!==a2));
  assign y11 = ((+(^(&$signed((!(~&(a1^b3)))))))!==(((b5&b4)>>(-a2))===$unsigned({b5,b5,a1})));
  assign y12 = ((a4?a2:a2)?(b1%a0):(a5?b1:p17));
  assign y13 = {3{p5}};
  assign y14 = {3{($unsigned((&(-{4{a3}}))))}};
  assign y15 = (3'd1);
  assign y16 = {(a4?a0:b0),(b3&&b4),(b5===a5)};
  assign y17 = (2'd3);
endmodule
