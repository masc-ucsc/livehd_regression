module expression_00162(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^(~&(3'd6)))?(&((4'sd5)^~(2'd2))):((4'd5)|(-4'sd4)));
  localparam [4:0] p1 = {3{{2{(-5'sd12)}}}};
  localparam [5:0] p2 = ((5'sd12)?{(4'd11),(-4'sd0),(-3'sd3)}:((3'd0)?(4'sd2):(5'sd2)));
  localparam signed [3:0] p3 = {((3'd5)^~(6'd2 * (2'd2))),(((3'd4)>>(5'd17))?(4'sd0):((3'sd2)^(3'sd3)))};
  localparam signed [4:0] p4 = ({((4'd13)!=(4'sd7))}>>>{(5'd2),(2'd2),(4'd12)});
  localparam signed [5:0] p5 = (((4'd12)<<<(3'd6))&((2'sd1)&&(4'sd4)));
  localparam [3:0] p6 = (-(5'sd2));
  localparam [4:0] p7 = (~&(~|{{2{{(2'd1),(-4'sd5)}}},{1{(~&(&(2'd2)))}}}));
  localparam [5:0] p8 = ((((2'd0)!=(4'd8))?((5'sd2)?(4'd0):(3'd1)):((-4'sd4)<(-4'sd4)))<<(((2'd1)&(-4'sd2))^((-2'sd1)!=(3'd6))));
  localparam signed [3:0] p9 = {(((2'd3)?(-3'sd2):(4'd5))===((3'd6)?(4'sd6):(5'sd8))),{{(2'd3),(4'd11),(2'sd0)}},(((2'd2)<=(2'd1))>{(-4'sd0),(3'd0),(3'sd0)})};
  localparam signed [4:0] p10 = ((((-2'sd0)^(5'd5))<(~(-(4'd7))))|(((5'd0)<=(3'sd1))?((4'd9)|(2'sd1)):((2'sd0)^~(-4'sd4))));
  localparam signed [5:0] p11 = (4'sd6);
  localparam [3:0] p12 = (-4'sd5);
  localparam [4:0] p13 = {(5'd22),{3{((4'd10)>>>(-5'sd10))}}};
  localparam [5:0] p14 = (((2'd0)>>>(-5'sd11))<{4{(2'd3)}});
  localparam signed [3:0] p15 = ((-5'sd6)&&(~^(~|((4'd11)&&(-3'sd1)))));
  localparam signed [4:0] p16 = {2{{{(5'sd3),(3'd1)},{1{(-4'sd5)}}}}};
  localparam signed [5:0] p17 = (~&(2'd3));

  assign y0 = {(4'd11),(5'sd1)};
  assign y1 = ($unsigned({4{p5}})<<$unsigned($unsigned(p11)));
  assign y2 = (3'd6);
  assign y3 = {{4{{a2,a1}}},(((4'd2 * a1)!=(p3<<b0))>>>({p4,a0,b1}+(b2<<b0)))};
  assign y4 = {2{{2{p12}}}};
  assign y5 = (&p10);
  assign y6 = ((((a0^p13)^(a0-p13))<{p8,p12,p4})<<<({(p15<<p13)}!=((p15&&b1)^~(b3!==b0))));
  assign y7 = (((4'd2 * b1)-{b2})>(~|(a4<p13)));
  assign y8 = {{1{((a5>>>b1)?{1{(3'd6)}}:(b0?a1:a2))}}};
  assign y9 = ($unsigned(((p12<=a4)+(p15!=b1)))>=$signed(({$signed((b2)),$signed((p4>p8))})));
  assign y10 = {(~|(~^(3'd7)))};
  assign y11 = ((((~a5)===(b1>>>b5))>{1{({4{b3}}>>>(a2<a5))}})==(|(~&(((b1<<<a0)&&{3{a2}})!==(+(b0<<a3))))));
  assign y12 = $unsigned($unsigned((2'd1)));
  assign y13 = {(|((~{2{p0}})>>>(2'd3))),((~&{{(p3>p17)}})|(|((&b1)>>(2'sd0))))};
  assign y14 = ((({p2,b3}?{1{b0}}:(p8+b5))|(&(p4?b3:p7)))>>(((~|p3)?(b2<<<b2):{p14,b0,p11})&&(~|((~&p10)>>>(~|p13)))));
  assign y15 = (p4?p14:p17);
  assign y16 = ({4{a1}}<<<(p1?b0:b0));
  assign y17 = (((|p13)<<<{4{b2}})?((|p11)!={4{p14}}):((!a1)||{3{p9}}));
endmodule
