module expression_00372(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'sd4)?(2'sd1):(4'd7))==={(~&(3'sd2)),((4'd4)?(4'd1):(2'd3))});
  localparam [4:0] p1 = {1{(5'd10)}};
  localparam [5:0] p2 = (((-2'sd1)?(2'd0):(4'd6))?((5'd17)?(5'sd4):(3'd0)):((2'sd0)?(-3'sd3):(5'd12)));
  localparam signed [3:0] p3 = (4'd13);
  localparam signed [4:0] p4 = (((5'd13)?(-4'sd2):(3'sd1))&((4'sd1)?(-2'sd1):(-2'sd1)));
  localparam signed [5:0] p5 = (+(((3'd1)<=(-5'sd6))<<((4'sd3)>(4'd9))));
  localparam [3:0] p6 = (((5'sd7)||(2'sd0))/(-5'sd5));
  localparam [4:0] p7 = ((-4'sd6)-(2'd2));
  localparam [5:0] p8 = {(2'd0),(5'sd14)};
  localparam signed [3:0] p9 = ((4'sd1)!=(5'sd8));
  localparam signed [4:0] p10 = (3'd3);
  localparam signed [5:0] p11 = (6'd2 * ((4'd8)^~(2'd0)));
  localparam [3:0] p12 = ((((3'd0)===(4'sd0))===(|(3'd5)))!==(5'd28));
  localparam [4:0] p13 = ((^((5'd28)%(-4'sd4)))>=((3'd0)>>>(5'd1)));
  localparam [5:0] p14 = (((-3'sd0)?(3'd1):(5'd25))?((4'd9)?(3'd3):(5'd4)):{4{(-5'sd4)}});
  localparam signed [3:0] p15 = (~^(~&({1{(((4'd0)>>(5'd27))|{4{(2'd0)}})}}<(((2'sd1)^~(-2'sd1))||{3{(4'd10)}}))));
  localparam signed [4:0] p16 = (-((^(+((3'd5)?(2'd3):(3'sd0))))<<(4'd7)));
  localparam signed [5:0] p17 = ((5'd13)===(3'd6));

  assign y0 = $signed(($signed($signed((|(a5==p3))))|((!p1)==(a4/b2))));
  assign y1 = (2'd1);
  assign y2 = (p17||p16);
  assign y3 = ((p7!=p10)>{4{p11}});
  assign y4 = {3{(^(-p16))}};
  assign y5 = {2{{{(3'd6)}}}};
  assign y6 = (|{4{(p12>b2)}});
  assign y7 = $signed($signed($signed((4'd6))));
  assign y8 = {{((p17^p2)<<{b5}),(-{3{p9}})},{{1{{4{b0}}}},{(!(b5||b2))}}};
  assign y9 = (|{4{((~^a3)<<(-a5))}});
  assign y10 = (!(-(&((6'd2 * (+(3'd1)))&&{(4'd9)}))));
  assign y11 = ((^((p13?p5:p12)?(p11?p4:p14):(a0?p6:a4)))||((5'd2 * p14)?(p11+p6):(p15^~p9)));
  assign y12 = $unsigned({1{{4{((p0?p2:b2))}}}});
  assign y13 = ((~|(~&{2{{1{b2}}}}))-(-((~|{2{p14}})<=(+(^b1)))));
  assign y14 = (&{((+(((b3?p15:a4))>{3{a3}}))+{3{{2{p16}}}})});
  assign y15 = ((p16<=p2)&(p5|p9));
  assign y16 = {(&(-5'sd7))};
  assign y17 = (p5<b3);
endmodule
