module expression_00889(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'd2)>>>(-5'sd7))=={(3'd0),(5'd0),(4'sd5)});
  localparam [4:0] p1 = (5'sd15);
  localparam [5:0] p2 = ((-4'sd7)>>(3'd7));
  localparam signed [3:0] p3 = ((2'd1)<<<(((-3'sd2)>>>(-4'sd1))!==((3'd5)<=(5'd23))));
  localparam signed [4:0] p4 = (&(((&((2'd0)^(2'd3)))>=(-(~&(2'd1))))<<<{2{((2'd0)<=(-5'sd4))}}));
  localparam signed [5:0] p5 = ((((3'd1)<<(4'd2))?(~^(5'sd15)):((4'd1)?(4'd14):(-4'sd0)))>=((&((5'd24)<=(5'sd10)))+((5'd12)?(5'sd1):(-5'sd13))));
  localparam [3:0] p6 = (2'sd0);
  localparam [4:0] p7 = ((2'd0)+(2'sd0));
  localparam [5:0] p8 = ({3{{(5'sd15),(3'd0),(5'sd5)}}}<<<((5'sd9)^~((3'd3)>(2'd1))));
  localparam signed [3:0] p9 = {4{((3'sd0)<=(3'd5))}};
  localparam signed [4:0] p10 = (+{1{({((4'd7)^~(3'd7)),(~&(4'd1))}-((4'd2 * (2'd0))||{3{(3'd0)}}))}});
  localparam signed [5:0] p11 = ((3'sd1)+(+((~^(-2'sd0))?((3'd2)?(4'd6):(3'd0)):((3'd2)^~(2'd2)))));
  localparam [3:0] p12 = (2'd1);
  localparam [4:0] p13 = ((((3'sd0)/(5'sd3))?((-3'sd3)?(2'sd1):(3'd3)):((2'd1)?(5'sd2):(-4'sd2)))?(((3'd3)-(4'sd6))?(&(4'sd4)):(|(2'd3))):(~(((5'd22)?(4'sd7):(5'd16))%(-3'sd2))));
  localparam [5:0] p14 = ((~|(~((4'sd2)==(-2'sd1))))&{{(-2'sd0),(4'd13),(-2'sd0)},((4'sd4)||(5'sd1))});
  localparam signed [3:0] p15 = ((~|{(-2'sd0),(-3'sd3)})|((~^(3'd3))>((-2'sd0)==(-3'sd2))));
  localparam signed [4:0] p16 = (({1{((-2'sd0)===(-3'sd1))}}<{4{(4'd14)}})^(((-4'sd3)+(-4'sd0))^((-3'sd0)?(4'd1):(3'd4))));
  localparam signed [5:0] p17 = (~^{{{{1{(-3'sd2)}}}},(-((-2'sd1)?(3'd3):(4'sd0))),(((3'sd2)?(5'd31):(4'sd2))<=((4'd12)?(3'sd3):(2'd0)))});

  assign y0 = (((b4<a4))!==($signed(b1)||(a0|a3)));
  assign y1 = ((~&(+p17))|((|p7)));
  assign y2 = (+$signed((-5'sd11)));
  assign y3 = ((~|(~^(~|(!(&p3)))))?(-({2{p9}}?(p17&p16):(p12||b3))):(-(+(p3?p5:p7))));
  assign y4 = (((3'sd2)+(a0>>p7))+$unsigned(((~|p11)<<<{4{b0}})));
  assign y5 = ((3'd5)==={(3'sd1),(2'd3)});
  assign y6 = (5'd30);
  assign y7 = (&(~(-(~|{4{(4'd10)}}))));
  assign y8 = ((b2?p2:p4)?(p0&p14):(~|(a1?p8:p17)));
  assign y9 = (((b2<<a2)?(b1&a5):(a5?a3:b4))==={4{(a5<a0)}});
  assign y10 = (-(((&p1)+(b4===a0))||($signed(a3)!==(~|b0))));
  assign y11 = ((b0<=b1)===(a5+b1));
  assign y12 = (((b5&&a2)!==(a1?b4:a5))?((p17<p10)||(a4+p11)):((p5?p6:p0)&(p16|p15)));
  assign y13 = {4{{(p9>>p17),(p2>>>p7)}}};
  assign y14 = {{({3{a1}}!==((a5<b0)<<(-5'sd2))),(-3'sd0)}};
  assign y15 = $signed($signed(((5'd2 * {2{a1}})+((4'sd4)==(p4)))));
  assign y16 = {(&{p4,p15,p6}),{1{(a3>p6)}}};
  assign y17 = {2{(p12?b1:b0)}};
endmodule
