module expression_00721(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((4'sd3)?(4'sd4):(2'sd1))};
  localparam [4:0] p1 = ((&((-3'sd1)>>(2'd0)))?((5'sd9)?(-4'sd0):(-4'sd5)):{2{(~(4'sd4))}});
  localparam [5:0] p2 = {{(4'sd7)},(5'd2 * (4'd6))};
  localparam signed [3:0] p3 = {3{(5'd5)}};
  localparam signed [4:0] p4 = ({2{((5'sd8)<(-4'sd1))}}<<<{{4{(3'sd0)}},{4{(4'd10)}}});
  localparam signed [5:0] p5 = (-(4'd11));
  localparam [3:0] p6 = ({{(5'sd4),(2'd2),(2'd2)},{(3'd3),(2'd1),(-5'sd4)}}==({(3'd5)}>>{(5'd18)}));
  localparam [4:0] p7 = ((~&({1{(5'd4)}}===((5'd25)^~(-5'sd4))))>(~^((-5'sd8)&(!(5'd12)))));
  localparam [5:0] p8 = {((((3'd2)^(5'sd3))!=((3'd6)?(4'sd2):(2'd0)))<<<(-2'sd0))};
  localparam signed [3:0] p9 = ((4'd15)-(2'd2));
  localparam signed [4:0] p10 = (4'd3);
  localparam signed [5:0] p11 = {1{(&{1{{2{(+((3'd7)?(-5'sd0):(-2'sd1)))}}}})}};
  localparam [3:0] p12 = ((4'd2 * {2{(5'd7)}})+{2{((4'd14)+(-2'sd1))}});
  localparam [4:0] p13 = (^(({(2'd2),(2'd3),(5'sd1)}+(-(+(3'sd0))))^(|(((-4'sd6)!==(-2'sd0))>=((4'd15)+(4'd5))))));
  localparam [5:0] p14 = {3{{(!((5'd20)-(-3'sd1)))}}};
  localparam signed [3:0] p15 = {{{{2{(5'sd9)}}}},(((5'd22)<<<(3'd4))<={(4'sd5),(-3'sd1),(5'd20)}),((-3'sd2)>>((3'sd1)>(2'sd0)))};
  localparam signed [4:0] p16 = (-(|(-(~&{((5'sd0)^~(3'd4)),{(5'd29),(-3'sd3)}}))));
  localparam signed [5:0] p17 = ((+{(3'd3),(2'd0)})===(-((2'sd1)&&(2'sd1))));

  assign y0 = {(3'd3)};
  assign y1 = (-$unsigned((&(5'd27))));
  assign y2 = (p14?p16:p8);
  assign y3 = (((b4?b1:b1)?(b0?b4:b3):(b0===a0))>=((a5)!==(~b1)));
  assign y4 = (~^({(&p14),(~&b0),{b1,p5,p0}}<<<{(b4||p6),(|a5),(p6<b4)}));
  assign y5 = {((6'd2 * (b1!==a1))^(+((3'd5)<<(4'd2 * p2))))};
  assign y6 = {1{{(~^p12),(-5'sd14),(3'd5)}}};
  assign y7 = {2{p8}};
  assign y8 = (~|(|(&((-(((p4))>(b3>>p3)))<=((~|(~&(-p3)))<<(&$unsigned((p11==p9))))))));
  assign y9 = ({p11,p6,a4}!=(~p8));
  assign y10 = (a2!=a0);
  assign y11 = ({{b3,p4,b4}}?(b3?p1:p5):(5'd2));
  assign y12 = (~{3{(b1?p15:p1)}});
  assign y13 = (4'd2);
  assign y14 = (~((p14&&p9)%a1));
  assign y15 = ({2{(a3<<p5)}});
  assign y16 = (5'd2 * {p6,p12});
  assign y17 = (-((b3|b0)==={2{b2}}));
endmodule
