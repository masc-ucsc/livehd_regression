module expression_00393(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(+((|(((5'sd1)|(4'd7))!=(5'd2 * (4'd12))))<<((4'd2 * (5'd4))>=(|(2'sd1))))));
  localparam [4:0] p1 = {((-4'sd5)<<(4'sd6)),((-3'sd0)<(4'sd5))};
  localparam [5:0] p2 = (~|((((2'sd1)<<(2'd0))-(~|(-4'sd7)))-((-4'sd2)||((2'd1)&&(-3'sd1)))));
  localparam signed [3:0] p3 = ((~{2{((3'd1)?(3'd1):(-3'sd0))}})?({(5'd24),(2'sd0)}&&{1{(5'd29)}}):{((2'd0)-(5'd19)),{(-4'sd2),(2'sd1),(3'd3)},((5'd20)!==(-3'sd0))});
  localparam signed [4:0] p4 = (+(2'd3));
  localparam signed [5:0] p5 = ((~(-3'sd3))?((2'd3)>>(5'sd10)):{(2'sd1),(4'sd7)});
  localparam [3:0] p6 = {2{(((5'd0)==(3'd7))!=={1{(-3'sd1)}})}};
  localparam [4:0] p7 = (((3'sd2)?(4'd0):(5'd23))^~((2'd2)<<(~(-3'sd3))));
  localparam [5:0] p8 = {(~&(5'd21)),((3'd7)===(5'd12))};
  localparam signed [3:0] p9 = ((!(2'sd1))<=(|(~^{(3'sd3),(3'd4),(4'd14)})));
  localparam signed [4:0] p10 = {1{{1{(3'sd1)}}}};
  localparam signed [5:0] p11 = ((((-5'sd15)<<(2'd1))<<((5'd8)-(4'sd2)))|(((-5'sd15)||(3'd2))!==((2'd0)>=(4'd8))));
  localparam [3:0] p12 = (~^((~(~((3'd6)<<<(5'd22))))!==(^(((3'sd1)<<<(2'd1))<<<((3'd1)-(5'sd12))))));
  localparam [4:0] p13 = {(2'd2)};
  localparam [5:0] p14 = (3'd1);
  localparam signed [3:0] p15 = {(({(3'd4),(2'd1)}||(~&(3'd6)))<<<((+(5'sd4))&&(~|(-4'sd4))))};
  localparam signed [4:0] p16 = (((-5'sd2)==(5'd11))>=((5'd21)^~(3'd7)));
  localparam signed [5:0] p17 = ((2'd3)|(5'sd3));

  assign y0 = ((~^b4));
  assign y1 = ({(~^{2{(p10==p9)}})}<<<(~&(~^(^{(p12>>p14)}))));
  assign y2 = (((a0===a1)?(p3<=p15):{p5})&((p9?p6:a4)?{b3,b2,p0}:(b3==a0)));
  assign y3 = $signed(a0);
  assign y4 = ($signed((-4'sd5))?((p16?a2:a4)?(p4?p10:b0):(-2'sd1)):(((-5'sd4)&(b3?p3:p6))));
  assign y5 = (~^((!(((!a3)&(^a1))-(^(p17>a1))))<(&((~&(a0>>>b1))>>(-(~(p17^~p4)))))));
  assign y6 = {(-4'sd0),{(5'd1),{a3,a0,a4}},(~&{{a4,a0}})};
  assign y7 = (~^(((b5==b4)<<<(b4<<a0))&((~^a3)-(~^a1))));
  assign y8 = ($unsigned({p5,p14,b4})?(5'd10):$unsigned((^$signed((p1)))));
  assign y9 = (~(|$unsigned(($signed(p3)))));
  assign y10 = ((((5'd2 * p8))|(p10&p15))&((p1|b5)>=(p11>>>p16)));
  assign y11 = {4{({4{p17}}?{1{p12}}:(b4?p14:p14))}};
  assign y12 = {2{a3}};
  assign y13 = {1{({2{(^{3{(~p17)}})}})}};
  assign y14 = (~(~^(((&$unsigned(p0))&&(b1<=b4))^~{(p15),(b0&&p12),(~^p12)})));
  assign y15 = $signed($signed((!((~|(-4'sd5))))));
  assign y16 = (2'sd1);
  assign y17 = ({2{(6'd2 * (!b2))}}>>>((~|(p3))?(a2^p5):(4'd2 * b2)));
endmodule
