module expression_00917(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd5)^~(2'd3))^((-5'sd14)?(2'sd0):(-2'sd1)));
  localparam [4:0] p1 = ({4{(2'sd1)}}>((-3'sd1)^~(-4'sd5)));
  localparam [5:0] p2 = (((-3'sd1)<=(4'd8))>>((-2'sd0)<<(5'sd13)));
  localparam signed [3:0] p3 = (((-5'sd12)^~(4'd3))<((3'sd1)!==(5'd27)));
  localparam signed [4:0] p4 = ((5'd2 * (4'd3))!==((2'd2)!=(-5'sd12)));
  localparam signed [5:0] p5 = (((-3'sd0)>>>(-5'sd15))^~(|(5'd1)));
  localparam [3:0] p6 = ((+(4'd13))?((-5'sd2)?(5'd8):(2'd2)):{{(4'd7),(5'd27),(4'd8)},(+(4'sd3))});
  localparam [4:0] p7 = (~&{1{{3{(5'd29)}}}});
  localparam [5:0] p8 = {({{(3'd0),(4'd5)}}<(&((4'sd1)>(5'd9)))),{{(-5'sd15),(2'd3),(2'd2)},{(4'd12),(-4'sd3),(4'd15)},{(5'd0),(5'sd8),(2'd1)}}};
  localparam signed [3:0] p9 = (~^(|(~(~|(~^(~^(~&(-(~^(~^(!(~^(-(~(2'd0)))))))))))))));
  localparam signed [4:0] p10 = (-(((3'd6)<=(3'd5))|(~^(3'd4))));
  localparam signed [5:0] p11 = (((2'd3)?(4'd1):(-3'sd3))?(^(+(4'sd2))):((-2'sd1)+(-4'sd6)));
  localparam [3:0] p12 = {4{({(-3'sd3)}!==((-5'sd10)?(5'd10):(3'd3)))}};
  localparam [4:0] p13 = {{((5'd22)||(4'sd0)),(((-3'sd0)==(3'd4))=={(5'd19),(5'd14)})},{((-5'sd15)>>(4'd5)),{(4'sd1),(4'sd5),(2'sd0)},((4'sd7)^~(-3'sd2))}};
  localparam [5:0] p14 = {{2{(+(6'd2 * (~&(!(4'd6)))))}}};
  localparam signed [3:0] p15 = ((((2'sd1)===(3'sd0))===((4'd2)>>>(3'd4)))-(((-3'sd1)<<<(3'd6))>=((2'd3)%(2'sd1))));
  localparam signed [4:0] p16 = {{(-4'sd6)}};
  localparam signed [5:0] p17 = (((5'd8)?(2'd3):(5'sd15))!=(((4'd5)?(2'sd0):(2'd2))|{1{(-4'sd0)}}));

  assign y0 = (b3>>p2);
  assign y1 = ({2{(b1?b1:a0)}}===((a4?a0:b3)?{b5,b4}:{b2}));
  assign y2 = (2'd1);
  assign y3 = $signed({1{{3{b3}}}});
  assign y4 = $unsigned(({1{$signed({1{{1{{4{p8}}}}}})}}));
  assign y5 = {1{b4}};
  assign y6 = {((p1-p11)>>>(p2>>>p15))};
  assign y7 = {{(p14||p10)},{3{p2}}};
  assign y8 = (~&(^{4{p4}}));
  assign y9 = ((|(a1>=a5))<={1{(b1===b2)}});
  assign y10 = ((~$unsigned((4'sd7)))>>>(((5'd13)<<$unsigned((p2>=b0)))));
  assign y11 = (~&((a5>p12)/p11));
  assign y12 = (p11+p0);
  assign y13 = (+{(~&(+((2'd1)>>>(~&p2)))),(-4'sd2),((5'sd11)<<<(3'd3))});
  assign y14 = {4{((~|p16)-(p4&&p8))}};
  assign y15 = (4'd14);
  assign y16 = ({2{(-2'sd1)}}?((p10?a3:a1)):((^p2)<<(2'd2)));
  assign y17 = ((-5'sd10)>(((a3?p16:b0)>(p12>=b2))||((p8&a3)&(-4'sd5))));
endmodule
