module expression_00407(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~&((4'd12)<<<(-4'sd0)))&(^((2'd0)<<(5'd8))));
  localparam [4:0] p1 = ({((4'd1)-(3'sd3))}===((!(5'd24))!=(!(5'd31))));
  localparam [5:0] p2 = {2{((4'd14)?(2'd0):(3'd6))}};
  localparam signed [3:0] p3 = (((3'd0)!=(4'd15))+((-3'sd2)<<(3'd0)));
  localparam signed [4:0] p4 = (6'd2 * {(5'd0),(5'd23)});
  localparam signed [5:0] p5 = ((4'sd5)<=(5'sd5));
  localparam [3:0] p6 = ({{(-2'sd1)}}?((5'd4)?(-2'sd1):(3'd1)):((-4'sd6)?(4'd15):(3'd6)));
  localparam [4:0] p7 = (-5'sd0);
  localparam [5:0] p8 = (2'sd1);
  localparam signed [3:0] p9 = ((~|{4{(5'd14)}})||(3'd3));
  localparam signed [4:0] p10 = {(!(&(((~&(3'd4))?((2'd0)!==(-4'sd2)):(~(4'd5)))!=((5'd2 * (4'd1))-{((5'sd8)^~(-2'sd1))}))))};
  localparam signed [5:0] p11 = ((3'sd3)===(4'sd2));
  localparam [3:0] p12 = (((3'd1)==((-3'sd3)<(3'd3)))!={((-3'sd2)!==(2'd3)),{(5'sd0),(-4'sd5)}});
  localparam [4:0] p13 = ((5'd5)-(3'd1));
  localparam [5:0] p14 = ((-3'sd1)%(2'd3));
  localparam signed [3:0] p15 = (((-4'sd7)==(3'd3))|((3'sd2)%(5'd1)));
  localparam signed [4:0] p16 = (2'd3);
  localparam signed [5:0] p17 = {4{(((5'd25)||(4'd11))&&{(-3'sd3)})}};

  assign y0 = (&((~|(~^(p11>>p12)))==(!(+(a5!==a0)))));
  assign y1 = ($signed(p17)?(p10?p5:p7):(p14^a0));
  assign y2 = (^(((~|{2{p4}})|{3{b3}})<({3{p2}}+{4{b0}})));
  assign y3 = (^{4{((^a2)?(p16<<<b0):(-p9))}});
  assign y4 = {{(p13||b3)},(&(b0+p4)),(-4'sd0)};
  assign y5 = (~{b0,a5});
  assign y6 = (|(((p9?p16:p9)<<(-4'sd1))?((b1?a1:a0)==={a5,a2}):(-(-5'sd15))));
  assign y7 = $signed($signed(p8));
  assign y8 = (~(~^$signed((~^$unsigned((~&((-5'sd5)^~$unsigned(b4))))))));
  assign y9 = (-(|(-3'sd1)));
  assign y10 = (|((~^{1{$signed(((b3-a4)))}})+$unsigned((|({3{b5}}>>>{2{p3}})))));
  assign y11 = (b2?b4:p12);
  assign y12 = {({p9,p0}<={p0,p17,p8})};
  assign y13 = (($signed((a5>>>b0))!==((~|b5)|(a1&a4)))!==((3'd0)));
  assign y14 = ((p8?p10:p8)|(p7+p12));
  assign y15 = (!(((p2^~a2)<(~b1))?((a1?a2:a5)>(b4>p15)):(&(b3?b5:b2))));
  assign y16 = (5'd17);
  assign y17 = (^(!(^((p17|p7)*(p5%a4)))));
endmodule
