module expression_00736(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(((4'sd7)>>>(4'sd6))<<<(^(2'sd0))));
  localparam [4:0] p1 = {4{{(-3'sd3),(-4'sd3),(5'd5)}}};
  localparam [5:0] p2 = (~&((^(~^(&(!(5'd11)))))==(~(((-2'sd1)&&(-5'sd7))&&{3{(4'd5)}}))));
  localparam signed [3:0] p3 = ((2'd1)<<((3'd4)?(-3'sd3):(4'd8)));
  localparam signed [4:0] p4 = ({4{(!(-3'sd3))}}&(({(2'sd0),(3'd2),(5'd23)}<={1{(4'd4)}})&&{(5'sd5),(-5'sd10),(4'sd7)}));
  localparam signed [5:0] p5 = ((-4'sd2)?{2{(4'sd2)}}:{4{(2'sd1)}});
  localparam [3:0] p6 = (~^{(~|(|({((4'd15)&(5'd2))}?((3'sd1)<<<(5'd11)):(-((5'sd9)&(4'sd7))))))});
  localparam [4:0] p7 = (-4'sd5);
  localparam [5:0] p8 = (+(+(-(+(~(-4'sd4))))));
  localparam signed [3:0] p9 = (((5'd2)|(-2'sd1))%(2'd1));
  localparam signed [4:0] p10 = (((-4'sd5)>=(-5'sd12))?{4{(-4'sd0)}}:(-3'sd2));
  localparam signed [5:0] p11 = ((+(-2'sd1))<<((2'd1)?(4'd6):(-4'sd6)));
  localparam [3:0] p12 = ((5'sd4)&(3'd0));
  localparam [4:0] p13 = ((-3'sd1)===((~((5'sd2)^~(5'd24)))<<<((4'd3)?(3'd5):(3'd1))));
  localparam [5:0] p14 = {4{(-5'sd3)}};
  localparam signed [3:0] p15 = (-((-4'sd3)<<(!(~|(-((!(2'sd1))<<<(4'd9)))))));
  localparam signed [4:0] p16 = {(!(3'd1)),((5'd18)!==(3'sd1))};
  localparam signed [5:0] p17 = {3{(((4'd13)?(-2'sd0):(3'd3))>=(&(4'd4)))}};

  assign y0 = ((5'd2 * (4'd2 * a1))>(((+(!a5))==={a0,b3})));
  assign y1 = ({2{{3{b4}}}}<(+{4{a4}}));
  assign y2 = $signed(p8);
  assign y3 = {(3'd5),{2{(-2'sd1)}},{3{(p17?b0:p2)}}};
  assign y4 = {(b5&a3),{p16,b4},{b4,a1}};
  assign y5 = {({b1,b3,a1}&(-4'sd7)),{{(p10<a3),(5'sd3)},{(b3?a5:b3),(b5<=p8)}}};
  assign y6 = {p3,p16,p6};
  assign y7 = ({1{$signed({4{{3{p13}}}})}});
  assign y8 = ((a3==a3)-$unsigned(a5));
  assign y9 = ({(~^(-2'sd1)),(|(b0?a3:a5))}-((-4'sd5)?(-5'sd11):(a1+b4)));
  assign y10 = ((-4'sd1)<<<(+{2{{2{p11}}}}));
  assign y11 = ((a5?a5:b0)<<<(5'd11));
  assign y12 = ((((4'd2 * p14))?(p3?a2:a5):$unsigned((p9<=p5)))<((p16^p16)?(p5>>>p17):((p17/p11))));
  assign y13 = {a2,b1};
  assign y14 = {(b5?b2:a1)};
  assign y15 = (({4{(a5?p8:p4)}}>>>((5'd11)&(b2+a4))));
  assign y16 = (2'sd1);
  assign y17 = (((b1!=a1)&&(a4!==a1))<<<{3{(5'd2 * p0)}});
endmodule
