module expression_00768(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(((-2'sd1)<<<(4'd4))!=((-2'sd1)!=(4'd14))));
  localparam [4:0] p1 = ((-{2{(+(5'd12))}})<={2{{4{(3'd0)}}}});
  localparam [5:0] p2 = ((|((4'd6)<<<(5'sd14)))^~((5'sd15)<(5'd0)));
  localparam signed [3:0] p3 = ((!((~&(-5'sd6))+((5'sd12)<(3'sd3))))>(4'sd4));
  localparam signed [4:0] p4 = ((5'd19)&(3'sd1));
  localparam signed [5:0] p5 = (+(~&(|(~|(~^(3'sd1))))));
  localparam [3:0] p6 = {4{{3{(3'd6)}}}};
  localparam [4:0] p7 = {2{({4{(3'sd0)}}?((2'd3)?(-5'sd6):(-5'sd10)):((-2'sd0)>>(4'd13)))}};
  localparam [5:0] p8 = (!((3'd1)^(((5'd30)&(3'sd0))?((5'd17)^(3'd7)):{(-5'sd11)})));
  localparam signed [3:0] p9 = {({(4'd0),(5'd1),(2'd1)}^~{((4'd9)+(-3'sd1)),{(2'd3)}}),((((2'sd0)^(4'd14))>>>((3'd7)===(2'sd0)))<((6'd2 * (2'd0))===((3'sd0)-(2'd3))))};
  localparam signed [4:0] p10 = (({1{((3'd5)>>(5'd10))}}+{1{{4{(5'd6)}}}})+{2{((-2'sd1)<<(5'sd3))}});
  localparam signed [5:0] p11 = {4{{1{((3'sd1)||(5'd4))}}}};
  localparam [3:0] p12 = ((((-4'sd4)&&(-2'sd1))>=((4'd5)<(-3'sd0)))<<((2'd2)?(4'd4):(-2'sd0)));
  localparam [4:0] p13 = ({1{{1{({4{(4'd5)}}>>>((4'd14)?(2'sd0):(-2'sd1)))}}}}<<<{4{((3'd7)>(2'd0))}});
  localparam [5:0] p14 = (+({3{(5'd23)}}!==(5'd2 * (5'd26))));
  localparam signed [3:0] p15 = ({3{(-4'sd4)}}?{4{(2'sd0)}}:((-2'sd0)?(-4'sd1):(4'sd4)));
  localparam signed [4:0] p16 = (~&((~|(((2'd0)>>>(4'sd2))?(~&(4'd11)):((4'd5)?(-3'sd2):(-5'sd4))))&&({(4'd15),(4'd14),(-3'sd1)}<((2'sd0)?(4'd1):(-3'sd2)))));
  localparam signed [5:0] p17 = ((|((5'sd12)<(-2'sd0)))-{1{{(2'd1),(-3'sd1)}}});

  assign y0 = (b3?a0:b0);
  assign y1 = ((~&(^(b1?p11:b4)))?(~&(~&(b3?b0:p5))):((-p3)?(&p6):{a2}));
  assign y2 = {{a3},(-b4),(~&a2)};
  assign y3 = {3{(3'd3)}};
  assign y4 = (a1>p2);
  assign y5 = {1{(3'd6)}};
  assign y6 = (((b0<=a4)^(+b0))>>>((a0*a0)>(a0|b3)));
  assign y7 = {4{(|$signed({3{b5}}))}};
  assign y8 = (5'sd12);
  assign y9 = ({{(p17?p14:b1),(a5?b4:p11),(~p0)}}?{(p12?p10:p11),(~^p9),{b3,p2}}:({b5,b4}^{p8,b1}));
  assign y10 = $unsigned($unsigned((+(|(~^$signed($unsigned((a0===b0))))))));
  assign y11 = ({{3{b2}},((+b2)),(a4?a0:b5)}===({3{a0}}?(b5?b0:b0):(|{b2,b1,b3})));
  assign y12 = {4{b1}};
  assign y13 = ((b2<<a5)<=(a4>a0));
  assign y14 = {2{((-$unsigned(b3))^~(a4>>>a3))}};
  assign y15 = (~^((4'd2 * (&{a1,b2,b2}))^~(((~|p10)!=(a0==b3))^~({(b2!==a5)}))));
  assign y16 = (4'd0);
  assign y17 = (&(|(5'd2)));
endmodule
