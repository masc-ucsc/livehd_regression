module expression_00300(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(2'd1));
  localparam [4:0] p1 = {4{((2'sd1)&&(-2'sd0))}};
  localparam [5:0] p2 = ((((-5'sd10)>>(-3'sd2))!=(3'd5))<<(-4'sd3));
  localparam signed [3:0] p3 = (|{{2{{(-4'sd0),(3'd2)}}},((+((4'd4)<<<(-2'sd0)))&{(^(5'sd0))})});
  localparam signed [4:0] p4 = {3{(~(|((5'sd0)>>(-4'sd0))))}};
  localparam signed [5:0] p5 = ((~&{2{((4'd11)?(3'd6):(-4'sd2))}})|(((2'sd0)?(3'd7):(4'd3))!=((3'd3)?(-5'sd0):(-5'sd15))));
  localparam [3:0] p6 = (({2{(5'd31)}}<{4{(-4'sd0)}})==(((-3'sd3)&&(2'd1))!=((-2'sd0)+(2'd0))));
  localparam [4:0] p7 = ({2{{(-2'sd0),(-3'sd1)}}}>({(-4'sd0),(4'sd0)}<={(4'sd3),(-2'sd1),(3'd0)}));
  localparam [5:0] p8 = ((6'd2 * (~|((3'd0)?(3'd0):(4'd2))))!=(!(2'sd0)));
  localparam signed [3:0] p9 = {3{(5'sd13)}};
  localparam signed [4:0] p10 = {(-4'sd3)};
  localparam signed [5:0] p11 = (((4'sd0)?(5'd9):(-4'sd2))?((3'd4)|(-2'sd1)):((3'd1)!==(3'd7)));
  localparam [3:0] p12 = {(4'd9),(5'd28)};
  localparam [4:0] p13 = ((|(~&((2'sd0)>>>(2'd0))))<<<({(4'sd3),(2'sd1)}|(~|(-2'sd1))));
  localparam [5:0] p14 = (5'd16);
  localparam signed [3:0] p15 = (2'd0);
  localparam signed [4:0] p16 = (~((^(-4'sd6))+(!(-(-5'sd0)))));
  localparam signed [5:0] p17 = (~&((-((3'sd0)==(3'sd1)))-((+(3'd2))^{1{(5'd23)}})));

  assign y0 = (~&(!(&(b4===b3))));
  assign y1 = (((4'd10)?(a4):(p5==b5))<<$signed(((b1?a1:a4)===(5'sd2))));
  assign y2 = ((2'sd0)?(4'd14):(~^(p11?a1:b0)));
  assign y3 = ((($signed($signed((p12>>a0)))==(-2'sd1))<=$unsigned((|(^((-b3)?(~&p5):(~^b1)))))));
  assign y4 = (~|$signed(({3{(^{4{p8}})}}|$unsigned({(~&$signed(b2)),(a4==p0),{2{p15}}}))));
  assign y5 = (({4{a3}}&(b4==b3))&(-2'sd0));
  assign y6 = {((5'd9)<((b0>>a1)!==(3'sd1)))};
  assign y7 = {$signed(((2'd1)>(~(5'd31)))),(-2'sd0)};
  assign y8 = (((4'd4)));
  assign y9 = ((!((b2?b2:a4)|(p14?p4:a1)))-((b3?b2:p15)?(~&b5):{3{p13}}));
  assign y10 = (((a4))!==$unsigned({b0}));
  assign y11 = (-4'sd5);
  assign y12 = $signed((-$unsigned({(!(|{3{p17}})),({3{a3}}),(^{$signed(b0)})})));
  assign y13 = (((p7<p14)?(a0?p16:b4):(b5?p0:p8))?((p4>a4)?(a2?p16:b0):(p4<<<p2)):((a4?a3:a5)==={4{a1}}));
  assign y14 = (3'd0);
  assign y15 = (~(!((p4+p1)>>>(-5'sd7))));
  assign y16 = {{b4,p10,p15}};
  assign y17 = (2'd1);
endmodule
