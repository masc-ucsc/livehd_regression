module expression_00456(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(-(~(2'd2)))}};
  localparam [4:0] p1 = ((2'd2)&{(-2'sd0),(5'd26),(2'sd0)});
  localparam [5:0] p2 = ((-((4'd12)>>>(2'sd1)))*((3'd7)<<<(3'd4)));
  localparam signed [3:0] p3 = (((-4'sd1)?(3'sd3):(5'd15))<<<(~^(2'd1)));
  localparam signed [4:0] p4 = (4'sd2);
  localparam signed [5:0] p5 = (((~&(-2'sd1))?{(3'd4)}:((3'd7)+(2'd3)))?{{4{(2'd2)}},{2{(-2'sd0)}},((5'd2)>(-3'sd3))}:(~((3'd0)?(4'd11):(5'd17))));
  localparam [3:0] p6 = {2{{(|(4'sd2))}}};
  localparam [4:0] p7 = (((2'd2)>>(2'd2))&(&(5'sd5)));
  localparam [5:0] p8 = (({{(4'd5),(5'd4),(-3'sd2)}}&{1{{2{(4'sd4)}}}})<<<(&(^({(-2'sd0)}===((5'd8)+(3'sd1))))));
  localparam signed [3:0] p9 = (~&((2'd3)?(3'd2):(5'd9)));
  localparam signed [4:0] p10 = ((~^(4'sd0))&&(^(-4'sd0)));
  localparam signed [5:0] p11 = (&(~|(!{4{((2'd3)>>>(-5'sd8))}})));
  localparam [3:0] p12 = (~|({3{(&(5'd30))}}^{4{(3'd7)}}));
  localparam [4:0] p13 = ((((3'sd0)?(5'd19):(2'sd1))?(^(-4'sd4)):(~^(4'sd1)))===((4'd2 * (2'd2))?((2'd3)-(2'sd0)):((4'd15)?(5'sd10):(2'sd0))));
  localparam [5:0] p14 = ((((4'sd2)==(5'sd7))>={{2{(4'd11)}}})=={4{((-4'sd2)==(2'd3))}});
  localparam signed [3:0] p15 = {3{(~(!((3'd7)?(-2'sd0):(-5'sd11))))}};
  localparam signed [4:0] p16 = (-(((5'd16)===(5'd3))>>(((4'd4)>(5'sd9))<<(5'sd14))));
  localparam signed [5:0] p17 = (((3'sd3)||(2'sd0))-((2'd2)<<<(2'd1)));

  assign y0 = {({1{a4}}^{1{p1}}),{(b4-b1),$signed(b0),$signed(a4)},((b1!==a1)=={p1})};
  assign y1 = (4'd12);
  assign y2 = (p16);
  assign y3 = {3{b4}};
  assign y4 = {(!{(-5'sd4),(a2>b4)}),(5'd11),(~^{3{(5'd16)}})};
  assign y5 = (~{2{(5'd2 * (~^$unsigned(b4)))}});
  assign y6 = ((|(p2?p12:p2))<(a3?p10:b4));
  assign y7 = (5'd8);
  assign y8 = ((p12+p10)&{2{p6}});
  assign y9 = (~|((&(($signed(b1)!=(~&b3))<<$unsigned((b4<<<p15))))));
  assign y10 = (5'd16);
  assign y11 = ((~&({4{b0}}!==((b1!==a3)||{2{a1}})))||((~^(b1<<b5))===((|a0)>>>(a3+a3))));
  assign y12 = ((~b0));
  assign y13 = (((a1^p12)<=(p15||p14))|((p5!=p8)!={p12}));
  assign y14 = (-{3{(&{4{b4}})}});
  assign y15 = (({{p14,p6},(!p0),$unsigned(b0)})?((^p10)?(a3&b4):(p0?a0:b1)):(~|((~|p2)?$unsigned(p16):(a1<<a4))));
  assign y16 = (-(^((p13?p6:a2)<<(b1?p16:a4))));
  assign y17 = ((4'd2 * (p0^b1))|(4'd2 * (b2^p2)));
endmodule
