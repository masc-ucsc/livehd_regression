module expression_00865(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(5'sd4),(3'sd1)};
  localparam [4:0] p1 = ((6'd2 * {(4'd0),(5'd7),(4'd13)})>(((3'sd2)?(-2'sd1):(4'd2))&&((3'd2)^~(-5'sd1))));
  localparam [5:0] p2 = ((~&(-2'sd0))>{(5'd26)});
  localparam signed [3:0] p3 = ((((5'sd7)>>>(2'd1))>>(~(5'd13)))==(((5'd30)+(-2'sd0))?((-2'sd0)>>>(3'sd1)):((5'sd10)?(-5'sd6):(5'sd3))));
  localparam signed [4:0] p4 = {2{(5'sd3)}};
  localparam signed [5:0] p5 = (3'd7);
  localparam [3:0] p6 = ((-(2'sd0))?(~|(2'd2)):((2'd3)?(-4'sd5):(-2'sd0)));
  localparam [4:0] p7 = ((!(~^(4'd0)))?(4'd2 * (5'd27)):(~^((-2'sd1)+(3'sd3))));
  localparam [5:0] p8 = ((2'd2)^~(3'sd1));
  localparam signed [3:0] p9 = (2'd3);
  localparam signed [4:0] p10 = {4{(-5'sd2)}};
  localparam signed [5:0] p11 = (((4'd12)===(-4'sd2))?{(-4'sd5),(4'sd2),(2'd3)}:((5'd11)>=(5'sd1)));
  localparam [3:0] p12 = (((~^(&(-5'sd1)))!==(4'd2 * (4'd14)))>>>((4'd8)!=(^((4'd2)>=(4'd7)))));
  localparam [4:0] p13 = ({((2'sd1)===(-4'sd1)),((3'd6)>>>(2'd1))}>=(((-2'sd1)+(5'd26))|{(3'sd2)}));
  localparam [5:0] p14 = (((4'd1)^~(4'd1))%(5'sd11));
  localparam signed [3:0] p15 = ((2'sd1)!=={(-5'sd7),(5'sd2),(4'd5)});
  localparam signed [4:0] p16 = (4'd1);
  localparam signed [5:0] p17 = (5'sd2);

  assign y0 = {({2{(^b5)}}?(^(-(~&a3))):{4{a3}})};
  assign y1 = ($unsigned((~&$signed(((~a0)?(p7?b3:a2):{4{a5}}))))|({b0,p16,p4}||{1{(p4>b4)}}));
  assign y2 = (((-p0)?(|a1):(p14))>>(~&(~&(b1?b4:a5))));
  assign y3 = (-4'sd7);
  assign y4 = (~^(|(~&(^(!{((p6^b1)&&{a5,p4,a1})})))));
  assign y5 = $unsigned($signed($unsigned($unsigned(((^(p17-p11)))))));
  assign y6 = (~|((!(p7?p7:p4))?(5'sd13):((p2?p0:p13)>>(-3'sd1))));
  assign y7 = {{b5,b5,p15},(2'd3),(4'sd2)};
  assign y8 = {4{a1}};
  assign y9 = ($signed((~^$signed(((p9^p16)^{p2,p2}))))||{(&(^(!(-(p5)))))});
  assign y10 = (-2'sd0);
  assign y11 = (p17?p13:b1);
  assign y12 = ((5'sd0)<<(4'd2 * (a0>>p2)));
  assign y13 = (!(-5'sd7));
  assign y14 = (~((&(p11?p17:b3))?(b3?a1:a1):(|{4{a0}})));
  assign y15 = {(5'd24),{1{{4{$unsigned(a5)}}}},{{3{p4}},$signed($unsigned(p0))}};
  assign y16 = $unsigned((~&(b2>>>b0)));
  assign y17 = ((3'd0)?(2'd3):(a1?b0:b2));
endmodule
