module expression_00758(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd12)|(4'sd0));
  localparam [4:0] p1 = ((3'd5)?(2'd2):(5'sd6));
  localparam [5:0] p2 = ((3'd3)<=(-3'sd0));
  localparam signed [3:0] p3 = (((3'd7)?(-4'sd4):(5'd21))!=((4'd14)!==(2'd1)));
  localparam signed [4:0] p4 = (~|(^(2'd0)));
  localparam signed [5:0] p5 = ({(5'd31),(2'sd1),(4'd0)}&&{(-2'sd1),(4'd11),(5'd18)});
  localparam [3:0] p6 = (-5'sd7);
  localparam [4:0] p7 = (^{1{(((-5'sd14)?(-4'sd6):(2'd3))!=((3'd4)?(-4'sd2):(5'sd0)))}});
  localparam [5:0] p8 = ((((-5'sd14)<<(4'd5))!=((5'd18)>(-4'sd5)))<<<(((4'sd7)||(3'd0))<<((3'd6)<<(-4'sd0))));
  localparam signed [3:0] p9 = (&((^((3'd5)&&(-5'sd6)))!==(((-2'sd0)^~(-3'sd2))>((-4'sd0)^(3'd1)))));
  localparam signed [4:0] p10 = ({3{(4'sd2)}}?((4'd4)===(-3'sd1)):((5'd1)+(4'd4)));
  localparam signed [5:0] p11 = {((|(5'sd6))||((4'd1)<=(-4'sd1))),(&{(2'd1),(3'd5),(4'd8)}),{1{{{(5'd18),(4'sd6),(3'd3)},(4'd10)}}}};
  localparam [3:0] p12 = ({1{{3{(~&(3'd5))}}}}||(!((-((2'd0)!=(-3'sd0)))^~{2{(2'd0)}})));
  localparam [4:0] p13 = ({1{{4{(2'sd0)}}}}=={4{(-5'sd10)}});
  localparam [5:0] p14 = {{((-3'sd2)>>(2'sd1))},(!{(5'sd14),(-5'sd8)}),({(-2'sd0)}^((-4'sd4)<<(4'd1)))};
  localparam signed [3:0] p15 = (^{4{(!(2'sd0))}});
  localparam signed [4:0] p16 = ((5'sd11)<(-2'sd1));
  localparam signed [5:0] p17 = ((+(((5'd30)<<(4'd15))?((-2'sd1)?(4'sd6):(2'sd1)):((-5'sd4)>(2'd3))))^~((-(-4'sd7))?(~|(4'd11)):(5'd2 * (2'd0))));

  assign y0 = (b0?p3:b5);
  assign y1 = (((&(~|p11))<={1{(p6<p11)}})!=($unsigned((p11))>(p1?p1:p12)));
  assign y2 = $unsigned((-2'sd1));
  assign y3 = ((a0!==a4)>(b5?a5:b3));
  assign y4 = $signed(b5);
  assign y5 = {1{{1{((+((b2<b5)>>>(a0!=a3)))!==(5'sd0))}}}};
  assign y6 = ((a5?p13:p9)?(3'd6):(|(p13>=p15)));
  assign y7 = {2{{{2{(b2>b1)}},{1{((a5>>a0)==={a3})}}}}};
  assign y8 = (|(-(4'd0)));
  assign y9 = {(a3?p6:a3),(b4||p15),{1{p11}}};
  assign y10 = ((&(b3&&p12))^~(!(+(p8^p13))));
  assign y11 = ((p13<=a5)?(|a0):(2'sd1));
  assign y12 = ((~(p8<b5))==(-(a3==a1)));
  assign y13 = {3{b5}};
  assign y14 = ((a4>>b1)==={a5,b3,a0});
  assign y15 = (4'd2 * {2{p1}});
  assign y16 = (4'd10);
  assign y17 = (^((($signed({p5,a3,a1})^~{$signed(a5)}))>>>{1{{4{{p11}}}}}));
endmodule
