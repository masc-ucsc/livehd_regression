module expression_00404(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((3'sd0)<(2'd2)),{{(-5'sd1)}},(2'sd0)};
  localparam [4:0] p1 = (-(+{2{{{3{(4'd3)}}}}}));
  localparam [5:0] p2 = ((((4'd3)?(2'd3):(-5'sd4))>>>((4'd6)?(4'sd1):(5'd18)))&&{1{(~|{4{(-3'sd3)}})}});
  localparam signed [3:0] p3 = ({(3'd5),(5'd12)}|((2'd2)&&(3'd6)));
  localparam signed [4:0] p4 = ((5'd8)?(-2'sd1):(5'd31));
  localparam signed [5:0] p5 = (~((4'd4)?(3'sd0):((-3'sd0)?(4'd12):(-2'sd1))));
  localparam [3:0] p6 = {1{((((3'd7)<(5'sd13))+((2'd3)===(3'sd2)))===(+({4{(3'sd2)}}-(~&(-5'sd4)))))}};
  localparam [4:0] p7 = ((-5'sd1)>>(4'd2 * (4'd2)));
  localparam [5:0] p8 = {({2{((3'd1)?(5'd8):(5'sd11))}}?{4{(2'sd1)}}:(4'd10))};
  localparam signed [3:0] p9 = {(-4'sd1),(4'sd7),(5'd3)};
  localparam signed [4:0] p10 = ((((3'sd0)?(2'd3):(3'd7))?((3'sd3)?(5'd24):(-4'sd4)):(~|(5'sd6)))||((5'd12)==((4'd4)==(-3'sd3))));
  localparam signed [5:0] p11 = (~|((2'd0)?(2'd3):(2'd1)));
  localparam [3:0] p12 = (^(-3'sd3));
  localparam [4:0] p13 = ((+{4{(&(-3'sd3))}})===(((2'sd1)>>(4'd14))=={2{(-5'sd8)}}));
  localparam [5:0] p14 = (5'd7);
  localparam signed [3:0] p15 = {2{((|(-(4'd3)))>>>{2{(4'sd2)}})}};
  localparam signed [4:0] p16 = (~|{4{((3'd2)?(2'd0):(4'sd0))}});
  localparam signed [5:0] p17 = {1{({3{((-5'sd5)>(-3'sd2))}}!=(((4'd2)|(2'd3))?{4{(3'sd1)}}:{2{(4'd10)}}))}};

  assign y0 = (2'sd0);
  assign y1 = ((b1^~b4)%a3);
  assign y2 = ((((a2^~a3)+(p3/a5))<$signed(((a4==a0))))==(($unsigned($unsigned(b2))/b4)));
  assign y3 = {(4'sd4)};
  assign y4 = (((p9>a3)>=(b0===a0))<=({a3,b0,p9}^(p4>b0)));
  assign y5 = ($signed($unsigned((~^(^(^(p16))))))==(~(~((p16<=p10)?(p10^~p13):(5'd23)))));
  assign y6 = $unsigned((((p4>=p6)?(b4==b0):(p9?p16:p11))?((b5!=b1)>>>(p16?p10:a5)):((p17?p13:p0)^~$signed($unsigned(p12)))));
  assign y7 = {4{{4{p3}}}};
  assign y8 = {1{(5'd2 * {3{p0}})}};
  assign y9 = ((a1?a4:a0)&&(b2?a4:p5));
  assign y10 = (((~^(a1!==b4))-(!(6'd2 * p2)))|({1{$unsigned(p12)}}>{4{p1}}));
  assign y11 = (((^(|p8))<={3{p13}})^~((~&p15)?(p14>>a3):{2{p7}}));
  assign y12 = (((-3'sd3)+(4'sd6))|(|(b0*a5)));
  assign y13 = {2{{4{p9}}}};
  assign y14 = ((({(p12>p4)})>>($signed({(p11||p15)})))|$signed($unsigned({{p16,p16},{p7,p10,p7},$signed({1{p4}})})));
  assign y15 = ((!((~&(b3&b5))<<(p11?b3:b4)))^~{3{(!(b2?a5:p9))}});
  assign y16 = {((-{(~&p17)})<{a0,p8,b1}),((&(p17>>b2))?(p7?a5:p16):(a2!=p15))};
  assign y17 = (~|{(!(+(^(!{(a4===b2)}))))});
endmodule
