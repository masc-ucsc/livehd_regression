module expression_00773(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd1)?(3'sd0):(5'd28))>>>((5'd11)^(3'd0)))!=(((4'sd5)*(-3'sd2))|((5'd16)<<(3'sd2))));
  localparam [4:0] p1 = ((~(((3'sd0)-(2'd2))^(~^(-2'sd0))))!=(((3'd5)||(-5'sd6))?(-(3'd6)):((-5'sd13)<<(5'd21))));
  localparam [5:0] p2 = ((-5'sd15)===(3'd4));
  localparam signed [3:0] p3 = {{3{(!(-2'sd0))}},(~&(5'd17))};
  localparam signed [4:0] p4 = {4{((4'sd3)^(-5'sd1))}};
  localparam signed [5:0] p5 = {(|(2'sd1)),((-3'sd1)==(5'sd1))};
  localparam [3:0] p6 = (((2'd0)?(5'd12):(-3'sd3))?((5'd15)?(5'd16):(5'd27)):((3'd7)?(-4'sd0):(3'd6)));
  localparam [4:0] p7 = (!({2{{2{(-3'sd0)}}}}!==(+(~((-3'sd3)+(5'sd2))))));
  localparam [5:0] p8 = (!((~|(~^{(3'd5)}))^~(5'd6)));
  localparam signed [3:0] p9 = (((~(4'd5))^((-3'sd3)<(2'd0)))^({(4'sd5),(5'd4),(5'd9)}||(+(-2'sd1))));
  localparam signed [4:0] p10 = (~&((4'd0)<=(-4'sd4)));
  localparam signed [5:0] p11 = (^{2{{2{{2{(-4'sd4)}}}}}});
  localparam [3:0] p12 = ({4{(2'sd1)}}==(((-4'sd2)&&(2'd2))<{2{(-5'sd2)}}));
  localparam [4:0] p13 = (~&(((2'sd0)||(3'd2))?(~&(4'd9)):(~&(-(-4'sd5)))));
  localparam [5:0] p14 = {4{((5'd28)>(3'sd2))}};
  localparam signed [3:0] p15 = {3{(4'd3)}};
  localparam signed [4:0] p16 = (((4'sd5)<<<(5'sd8))%(4'd1));
  localparam signed [5:0] p17 = ((-3'sd3)?(5'sd6):{(4'd12)});

  assign y0 = {({p13,a0,p7}||(b0?p9:b1))};
  assign y1 = (p5?a5:b0);
  assign y2 = (5'd14);
  assign y3 = (~^((&(~|(~^(^p16))))^~(|(~&(p12>=p7)))));
  assign y4 = (|{p7,p5,a0});
  assign y5 = (3'd0);
  assign y6 = (((2'd3)>(a5>>b3))==={1{{1{(b0<b0)}}}});
  assign y7 = (((~^b5)?(4'sd1):(p11))>((2'd2)>=(b1||p4)));
  assign y8 = (^(~|a4));
  assign y9 = (($unsigned((a3*a1)))!==(2'sd1));
  assign y10 = $unsigned({$signed(((+(a1<=p14))+(a0?p9:a4)))});
  assign y11 = (((a5)!==$signed(b4))>$signed($unsigned((5'd2 * b0))));
  assign y12 = (($signed(b0)!=(b0?a0:a1))?$unsigned((a5^b5)):(p4?a2:a0));
  assign y13 = (~|(($unsigned((b3>>>p17)))?{((p15?p7:p17)<<(^a4))}:((~|a1)&(~^p13))));
  assign y14 = (|{2{(-2'sd0)}});
  assign y15 = (~|a0);
  assign y16 = {4{{3{{3{b0}}}}}};
  assign y17 = (~|a3);
endmodule
