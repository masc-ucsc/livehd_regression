module expression_00293(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd0)!==(5'd2))||((5'd20)-(2'd2)));
  localparam [4:0] p1 = (+(((~&(-2'sd1))?(~&(-5'sd14)):(4'd2 * (2'd2)))?((5'sd2)?((5'sd2)>=(-4'sd6)):(&(-2'sd0))):((4'd1)?(2'd3):(!(4'd4)))));
  localparam [5:0] p2 = ({2{{2{(5'd14)}}}}!==(((3'd2)?(5'd1):(3'd6))?((3'sd3)?(5'd19):(3'sd1)):{4{(3'sd1)}}));
  localparam signed [3:0] p3 = {{(3'sd2),(2'sd0)},((-3'sd1)?(2'd0):(2'sd0)),(!(2'd2))};
  localparam signed [4:0] p4 = {(4'd2 * ((3'd1)^(4'd1)))};
  localparam signed [5:0] p5 = (~|(5'd9));
  localparam [3:0] p6 = (4'd15);
  localparam [4:0] p7 = (-((-3'sd2)!=((5'd27)&(3'd0))));
  localparam [5:0] p8 = ((!((2'sd1)^~(-2'sd1)))!={3{(-2'sd1)}});
  localparam signed [3:0] p9 = (+(~{(&(~^{((&{3{(-5'sd11)}})-(~^(((2'd0)^~(5'd6))<<(~^(5'd4)))))}))}));
  localparam signed [4:0] p10 = {(3'd1),(-4'sd5),(4'sd5)};
  localparam signed [5:0] p11 = (|(~|((2'sd1)<<<{4{(5'sd0)}})));
  localparam [3:0] p12 = ((((2'd0)>>>(2'd2))|{1{(5'sd9)}})?(-4'sd4):({4{(5'sd8)}}?{(5'd16)}:((3'd3)?(-2'sd0):(5'sd2))));
  localparam [4:0] p13 = (+(~&(4'd7)));
  localparam [5:0] p14 = {({{(3'd7),(5'd1)},((2'd1)||(2'sd0)),{(2'd3),(5'd10),(4'sd3)}}===(((3'd3)+(3'sd1))^~((-5'sd0)>>(2'sd0))))};
  localparam signed [3:0] p15 = ((2'd1)<=(5'sd7));
  localparam signed [4:0] p16 = ((((-2'sd1)&(2'd1))<=(-3'sd1))>((-3'sd1)<<{(-5'sd5),(4'd0),(2'd1)}));
  localparam signed [5:0] p17 = (~(^(-2'sd0)));

  assign y0 = ((5'd13)<=({2{(~^a0)}}||(^(~&(p7?a4:p11)))));
  assign y1 = (3'd2);
  assign y2 = (^{(&{3{{3{(p5?p0:p0)}}}})});
  assign y3 = ({4{p6}}?(-p12):(~&p9));
  assign y4 = (((b1+p8)+{1{p2}})?((4'd2 * p13)):((&p12)>>(+b4)));
  assign y5 = (|((((4'd13))/p8)?(^(|(4'd11))):(~&(4'd5))));
  assign y6 = $unsigned((((p16|p3)?(~^p9):(p8!=a0))<<((&p7)?(p11?p4:p14):(p5-p17))));
  assign y7 = (((4'd2 * (a2|a1)))!=$unsigned(($signed($signed(p14))/b5)));
  assign y8 = {4{{1{{1{b3}}}}}};
  assign y9 = $signed(((3'sd2)));
  assign y10 = (|({4{b0}}!==((b0)===(a4>>>a2))));
  assign y11 = {2{((~^p16)>(b4!==b2))}};
  assign y12 = $signed(({($unsigned({3{p5}})<<<$unsigned((p2|p11)))}<(((a4!==b1)>=$signed(a4))>>(4'd2 * $unsigned(b3)))));
  assign y13 = (~((p1+p2)?(a4?p10:p16):(-3'sd1)));
  assign y14 = (({{3{p16}}}<={{p13,p5},(p9>p5)})>>(({2{p0}}>>{1{p6}})>={(5'd2 * p6),(p8&&p2),(b5!==a1)}));
  assign y15 = (~^((|(|(~|(+(2'd1)))))?(|$unsigned((-(-(|p5))))):({2{p2}}?(p9?a1:p14):{4{b3}})));
  assign y16 = ((|(|(a3>p10))));
  assign y17 = $unsigned($unsigned({((p11?p9:p6)?$signed(p6):(2'd1)),((p17>>p10)?(4'd6):(p10^~b4))}));
endmodule
