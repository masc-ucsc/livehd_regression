module expression_00894(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({4{(2'd2)}}&{(2'sd1),(2'd3),(4'sd5)})?{4{(5'sd13)}}:({(3'sd0)}?((-2'sd0)+(4'd15)):((4'd2)>(4'd5))));
  localparam [4:0] p1 = (((2'd1)?(-4'sd5):(-4'sd4))?((-3'sd1)?(3'd6):(4'd5)):(~^((-4'sd7)?(2'd2):(-5'sd15))));
  localparam [5:0] p2 = (((-4'sd0)>>(~&((4'sd1)<<<(-2'sd0))))===(4'd3));
  localparam signed [3:0] p3 = (((~&(4'sd7))!={2{(2'sd1)}})?(4'sd0):((-(2'd2))>=(!(4'sd3))));
  localparam signed [4:0] p4 = (~|(((5'd27)<(-5'sd11))?((-4'sd2)<(3'sd2)):((-3'sd1)>(2'd1))));
  localparam signed [5:0] p5 = (3'd1);
  localparam [3:0] p6 = {{{4{(-3'sd1)}},{(-3'sd1),(2'sd0),(-5'sd0)},({3{(2'd2)}}===((-3'sd3)^~(5'd8)))}};
  localparam [4:0] p7 = (!{1{(4'd12)}});
  localparam [5:0] p8 = (3'd3);
  localparam signed [3:0] p9 = {((2'd0)&&(!({(~(3'd3))}&(5'd10))))};
  localparam signed [4:0] p10 = ((3'd0)?((-4'sd5)?(-2'sd1):((-2'sd0)<<<(2'sd0))):{((-5'sd15)<(-5'sd2)),((3'd4)===(2'sd0))});
  localparam signed [5:0] p11 = (3'sd1);
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = (2'd1);
  localparam [5:0] p14 = (~&((-(((2'd2)>=(4'sd2))===((3'd1)^(3'sd1))))>>>(|(^((-2'sd0)+(4'd5))))));
  localparam signed [3:0] p15 = (((-2'sd0)<=(4'sd2))||{4{(4'sd0)}});
  localparam signed [4:0] p16 = {(-3'sd2),((-3'sd3)?(-5'sd15):(5'd4))};
  localparam signed [5:0] p17 = ((((-5'sd4)>>(-5'sd10))-((5'sd2)>>>(2'd1)))?{{(2'd1),(4'd0),(-4'sd3)}}:(((2'sd1)>=(2'sd0))?(6'd2 * (3'd7)):((5'd10)|(-2'sd0))));

  assign y0 = (~((~&({2{b4}}?{1{$unsigned(p3)}}:$signed($unsigned(b1))))==(~{3{(p5?p17:p8)}})));
  assign y1 = {4{(-{1{(a2===b5)}})}};
  assign y2 = ({(p8?p2:p13),(~p12),{p0,a3,p9}}?{4{(p17<<<p17)}}:{(&(4'sd3)),{p13,p3}});
  assign y3 = {3{(4'd2 * $unsigned($unsigned(a5)))}};
  assign y4 = (~|((~|(a0?a2:p10))-((|b4)>>>(p4?p12:p0))));
  assign y5 = (({p1,p7}<<<{p4})=={p3,p7,p14});
  assign y6 = {3{$unsigned(((p6)<={4{b2}}))}};
  assign y7 = (~&{4{(~$signed((!$signed(b5))))}});
  assign y8 = ((p2+p15)&&(p13>p3));
  assign y9 = {1{{3{((+{3{p8}})>=(&(5'd19)))}}}};
  assign y10 = {({2{b5}}!=({4{a1}})),((a4<<<b0)^~(b0^~b4))};
  assign y11 = (((b3?p8:p16)<<<(p15||p4))?(2'd0):((p11<=p2)?(-5'sd1):(b3-p8)));
  assign y12 = (p3<<<p12);
  assign y13 = (!((+((~(+a1))&&(~|(!a3))))==((b0/b3)%b2)));
  assign y14 = ((-{(((a2===b2)+(p4?b1:p6))&(p11?a4:p12))})^(6'd2 * (p6?p0:p7)));
  assign y15 = ((+(b3%p16))%b0);
  assign y16 = {3{((b5?p15:p9)?(b5?b3:p14):$unsigned(p13))}};
  assign y17 = (!({2{a0}}));
endmodule
