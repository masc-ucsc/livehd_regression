module expression_00409(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-4'sd0);
  localparam [4:0] p1 = (((-2'sd1)%(-3'sd2))?((-4'sd2)?(-3'sd3):(5'sd6)):((2'd3)!==(3'd0)));
  localparam [5:0] p2 = (({4{(-5'sd11)}}>>>(4'sd3))>>>{2{((4'sd5)^(2'sd0))}});
  localparam signed [3:0] p3 = (^(&(~^(~&(!((~&(!((-5'sd2)|(-3'sd0))))-((~^(-4'sd5))*(~^(2'sd0)))))))));
  localparam signed [4:0] p4 = ((-5'sd15)^(2'd2));
  localparam signed [5:0] p5 = ((!((5'd29)+(-4'sd2)))?{1{((5'd18)<<(-2'sd0))}}:{1{(&(^(4'd14)))}});
  localparam [3:0] p6 = ((^(!{((2'd0)?(5'd29):(2'd0))}))?((^(-4'sd5))>>{(-2'sd0),(5'd15),(3'd5)}):((&(-4'sd0))?((4'd10)?(3'sd2):(-2'sd1)):((4'd14)?(3'd4):(5'd28))));
  localparam [4:0] p7 = {((2'sd0)?(-2'sd0):(3'sd3)),{3{(3'd2)}},({2{(-5'sd2)}}||((2'd3)<<<(-2'sd0)))};
  localparam [5:0] p8 = (5'd17);
  localparam signed [3:0] p9 = {((~|(6'd2 * (5'd12)))&&{(3'sd2),(-5'sd12)}),{(((5'sd6)^(5'd19))<=((4'd4)<<<(-4'sd4)))}};
  localparam signed [4:0] p10 = (((-5'sd0)<<<(4'd14))+((-2'sd1)===(2'd0)));
  localparam signed [5:0] p11 = (-4'sd1);
  localparam [3:0] p12 = (((4'd13)<<<(-5'sd11))^~{(5'sd0),(5'd9)});
  localparam [4:0] p13 = {(~^({(5'd10)}^~((3'd5)>>(5'd16)))),(-(5'd2 * ((3'd1)&(3'd0))))};
  localparam [5:0] p14 = ((((2'd1)^~(-4'sd3))-((3'd3)<=(-4'sd5)))>>((-5'sd0)?(4'd15):(3'd3)));
  localparam signed [3:0] p15 = ({3{(2'sd1)}}>>((5'd5)<<(4'sd7)));
  localparam signed [4:0] p16 = (4'd6);
  localparam signed [5:0] p17 = (|(!(^(5'sd5))));

  assign y0 = {3{(-5'sd6)}};
  assign y1 = (-(p1&a3));
  assign y2 = {({b3,b4,b0}?(-3'sd1):(b4>p8)),{2{{a4,a0,a1}}},(-4'sd0)};
  assign y3 = {3{b1}};
  assign y4 = {3{(!p8)}};
  assign y5 = (b4?b4:b4);
  assign y6 = {({p6,a1,a4}<<(a2<<b3)),({a5}&(2'd3)),$signed((-(5'd22)))};
  assign y7 = {{{1{(p14?a2:p5)}},(p7?p5:a2)},((-5'sd10)!==((a1&a3)&(a5>b2)))};
  assign y8 = (3'd4);
  assign y9 = (3'd0);
  assign y10 = (4'd6);
  assign y11 = (((-2'sd0)?{a5,b2}:{b4,a5})-((3'sd1)));
  assign y12 = {2{(5'd22)}};
  assign y13 = (~^{(p8>>>a3),(p13?p5:p13)});
  assign y14 = (((p2<<<p0)>>>(a1?b4:a3))?{3{a1}}:{1{(-(~&a1))}});
  assign y15 = $signed((~&{1{{2{((b4===a1)<(p1?p12:p4))}}}}));
  assign y16 = ((|{b3})+(b2?p8:a0));
  assign y17 = ({(p17|p8),(p11?p12:p7)}>>{1{{4{p5}}}});
endmodule
