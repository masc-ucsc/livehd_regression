module expression_00459(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{(-3'sd3),(5'd17)}}};
  localparam [4:0] p1 = (-4'sd5);
  localparam [5:0] p2 = {{((4'd1)!={(-4'sd3),(3'sd1),(4'd3)}),(4'sd2)}};
  localparam signed [3:0] p3 = ((({(-2'sd1),(4'd3)}&&(5'd21))|{((3'd7)<<(4'sd0)),((-3'sd3)<<<(4'sd5))})&(((2'sd1)?(3'd1):(-4'sd2))?((-4'sd5)?(3'sd2):(3'sd0)):((5'sd7)<(-5'sd1))));
  localparam signed [4:0] p4 = {(3'd6),(5'd3),(3'sd0)};
  localparam signed [5:0] p5 = (6'd2 * ((5'd3)^~(5'd11)));
  localparam [3:0] p6 = {{{(-4'sd2),(2'd2),(4'd11)},{((-4'sd7)?(5'd13):(-4'sd3))},(~^(~&(-(-3'sd3))))}};
  localparam [4:0] p7 = (~^(+(^{4{{1{(&(5'd3))}}}})));
  localparam [5:0] p8 = ({1{(((5'd30)<<<(4'd1))===((2'd3)||(5'sd12)))}}<(((2'd3)>>>(4'd14))||{(-2'sd1),(2'd3),(5'sd13)}));
  localparam signed [3:0] p9 = (|(+((((-4'sd5)===(-4'sd2))>>>{1{{4{(4'd6)}}}})<{2{{3{(4'd13)}}}})));
  localparam signed [4:0] p10 = ((((4'd11)&&(-2'sd0))^((5'd27)<(-3'sd2)))||(((3'sd2)>(4'd14))*((4'sd2)&&(-5'sd9))));
  localparam signed [5:0] p11 = (((3'sd2)+(2'sd0))^~(-4'sd0));
  localparam [3:0] p12 = (3'd2);
  localparam [4:0] p13 = ({2{(4'd2 * (3'd5))}}+({1{((3'd1)<<(3'd3))}}<((2'sd1)!==(2'd3))));
  localparam [5:0] p14 = {2{{(5'sd5),(-5'sd1),(-2'sd0)}}};
  localparam signed [3:0] p15 = (((2'd0)%(2'd1))^~(3'd6));
  localparam signed [4:0] p16 = {((3'd7)<=(5'd1)),(^((-4'sd0)<(-4'sd4))),{2{(2'd3)}}};
  localparam signed [5:0] p17 = (|(5'd9));

  assign y0 = (((a0!==b4)!==$signed((4'sd5))));
  assign y1 = {(~|(!(!p8))),{((^p12))}};
  assign y2 = ((~({(a4+p3)}=={p13,p8,p11}))<=((a1===a1)+(p4<<p3)));
  assign y3 = (((!b0)>=(b0<<<b4))!==((-b5)<<<(a0*a5)));
  assign y4 = (^(!(&{4{(&b0)}})));
  assign y5 = ((b5>>>a0));
  assign y6 = (({1{p4}}<=(a5<<p7)));
  assign y7 = {(-2'sd0),({3{p7}}?{4{p11}}:{p12})};
  assign y8 = {2{((5'sd1)<<{3{a4}})}};
  assign y9 = (5'sd6);
  assign y10 = (6'd2 * $unsigned({p14,p6,p14}));
  assign y11 = (+(4'd4));
  assign y12 = (3'sd2);
  assign y13 = ({{p17,b3,p14}}==(b3^~p13));
  assign y14 = {{(~{2{(|(~&(^p16)))}})}};
  assign y15 = (~^{b2,b3});
  assign y16 = (p1-p0);
  assign y17 = $signed(($unsigned((((-4'sd6)<(b3?p8:p7))))?((3'd2)?(5'sd10):(5'sd11)):(3'd4)));
endmodule
