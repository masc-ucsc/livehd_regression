module expression_00160(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-{(4'd4),(-2'sd0),(4'd9)});
  localparam [4:0] p1 = (((5'sd4)<(3'sd3))>=((4'd3)>(2'd0)));
  localparam [5:0] p2 = ((4'sd1)?(4'sd4):(-4'sd7));
  localparam signed [3:0] p3 = (-4'sd6);
  localparam signed [4:0] p4 = ((~&{4{(5'sd0)}})?(!(((-5'sd7)>=(2'sd1))===((5'd11)?(3'sd1):(4'sd7)))):{2{((4'd4)!=(5'sd9))}});
  localparam signed [5:0] p5 = (2'd0);
  localparam [3:0] p6 = ((((4'd4)?(2'd1):(4'sd3))||{1{(-3'sd0)}})?(((5'd10)>=(-2'sd1))?((3'sd0)^~(-4'sd5)):((5'sd13)===(4'sd2))):({1{(4'sd3)}}?((4'd3)?(-4'sd3):(-4'sd1)):((5'sd7)>>(5'd14))));
  localparam [4:0] p7 = (2'd2);
  localparam [5:0] p8 = ((2'd3)<(-5'sd3));
  localparam signed [3:0] p9 = (({(4'd13),(5'd14),(3'sd3)}==((-5'sd7)>>>(2'd3)))<(((5'd15)!==(5'd12))+{(3'd4),(4'd4),(4'sd7)}));
  localparam signed [4:0] p10 = (-(+(((4'd14)?(3'd1):(2'sd0))*(&(+(4'sd4))))));
  localparam signed [5:0] p11 = (((6'd2 * (2'd0))+((4'd5)?(4'd1):(-3'sd2)))|{1{(&(^{1{(4'd2 * (2'd1))}}))}});
  localparam [3:0] p12 = (~&((((-3'sd3)<(5'sd14))^~((-2'sd1)<<(2'd2)))>=(((-3'sd1)&(5'sd5))<<<((-4'sd2)^(-2'sd0)))));
  localparam [4:0] p13 = ((|(((3'd7)<<<(2'd2))?((3'd7)+(-3'sd3)):((4'd15)<<<(-4'sd5))))-(((4'd7)?(-2'sd1):(-5'sd4))&&((3'd0)?(2'sd0):(3'sd0))));
  localparam [5:0] p14 = (3'd1);
  localparam signed [3:0] p15 = ((((5'd10)>(-4'sd1))&((2'd2)-(-5'sd5)))===(2'sd1));
  localparam signed [4:0] p16 = (2'd3);
  localparam signed [5:0] p17 = (|{3{((-5'sd9)?(-4'sd2):(-2'sd1))}});

  assign y0 = {4{((a2>=b1)^(~|b1))}};
  assign y1 = (-5'sd3);
  assign y2 = (3'sd1);
  assign y3 = (3'sd1);
  assign y4 = {2{{2{{2{(b2>=b5)}}}}}};
  assign y5 = ((((a4<<<b5)^(b4-a0))!==((a4^a2)^(+a0)))<<<(({p11}+(~^p5))&&((p7==p3)-(p11^p11))));
  assign y6 = $unsigned((({3{$signed(p15)}})));
  assign y7 = {(|(~&(~&({p14,p17}?(p8==p1):{a5,p2,p0})))),(~((p3?p17:p7)?(p16&p15):(~^(p6?p10:p9))))};
  assign y8 = {(-{((a0===b3)!=(!a0)),{(-(b0<<<p6))}}),((&(!(-(+a5))))>=(|({b2,b2,b2}|(a1==p7))))};
  assign y9 = (a4?a2:p0);
  assign y10 = (2'sd1);
  assign y11 = (((b1<<<a3)<<(b4>>>p0))?((b3?b5:b0)<<(b3===a4)):((a3==b4)>>(b3!=a3)));
  assign y12 = (|(+(((3'd7)))));
  assign y13 = {1{(!(&b1))}};
  assign y14 = ($unsigned(($unsigned({p17,a0,p0})?(p3?p0:p1):(p1^p17)))<<<{((p5?a0:p2)>=($signed(b2)^~(p14+b1)))});
  assign y15 = {p15,p12,p1};
  assign y16 = ((p13?p15:p5)<=(p6?p13:p7));
  assign y17 = ($signed({((p17)>>>(p0^a1))})<{{a4,p2,a2},{1{b0}},{p13,b4,p15}});
endmodule
