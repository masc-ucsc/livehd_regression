module expression_00329(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd1);
  localparam [4:0] p1 = (|(~(2'd1)));
  localparam [5:0] p2 = (^(3'd5));
  localparam signed [3:0] p3 = ((((2'd2)<=(-5'sd15))^~(~(4'd10)))<={{(3'd2)},((-2'sd1)+(3'd0))});
  localparam signed [4:0] p4 = (3'd0);
  localparam signed [5:0] p5 = ((^(4'd9))?((-4'sd0)&&(2'sd1)):((-3'sd1)&(2'd3)));
  localparam [3:0] p6 = ((5'sd14)<<<(~(~((4'd12)!=(-5'sd9)))));
  localparam [4:0] p7 = ((~&((5'd2 * (3'd5))|(~(5'd27))))<={(!(-2'sd0)),{(3'd1),(3'd7)},((2'd1)||(-3'sd2))});
  localparam [5:0] p8 = (({(4'd5),(4'sd0)}?(~|(-3'sd2)):((2'd3)==(5'd0)))>>>(((4'd14)<<<(3'd7))&((-2'sd0)>(4'sd4))));
  localparam signed [3:0] p9 = ({((3'd5)^~(5'd5)),((-4'sd3)+(2'sd1))}=={{{(2'd0),(5'd9),(-3'sd3)},((3'sd3)==(-2'sd0)),((2'd0)>>(4'sd4))}});
  localparam signed [4:0] p10 = (((-2'sd0)?(4'd12):(2'sd1))^((4'sd2)<<(4'sd1)));
  localparam signed [5:0] p11 = ({((3'd7)?(3'd0):(5'd26)),(-(-3'sd1))}?({(5'd15),(5'd19)}==((5'd11)&&(4'd13))):((~(3'sd2))<<<((5'sd3)===(4'd9))));
  localparam [3:0] p12 = ((({1{(3'd3)}}<{(5'sd10),(5'd10),(2'sd0)})>>({3{(2'sd0)}}<<<{2{(2'sd0)}}))>({(-{(5'sd8),(5'd25)})}>>>{3{(5'sd14)}}));
  localparam [4:0] p13 = ((~|(((3'sd2)==(5'd8))===((3'd0)>=(-2'sd1))))&(+(~|((5'd10)>(4'd11)))));
  localparam [5:0] p14 = ((|(((3'd3)===(-5'sd5))?((3'sd2)?(5'd2):(-2'sd0)):(|(3'sd1))))>={{(4'd10),(-3'sd0),(-2'sd1)},{(4'sd3)},(&(5'sd4))});
  localparam signed [3:0] p15 = (!{2{(!(4'd0))}});
  localparam signed [4:0] p16 = ((((4'd8)<<(4'd1))&((4'd3)^(-2'sd0)))>>(((-5'sd15)^(-2'sd1))>>((3'd3)%(4'd0))));
  localparam signed [5:0] p17 = {(2'd2),(2'sd1),(5'sd2)};

  assign y0 = {(+(2'd1)),{1{{((5'd28)?(a2==a5):(a4>>>b0))}}}};
  assign y1 = (((b4)-(p4?b5:p2)));
  assign y2 = (6'd2 * (~^(a2^~a2)));
  assign y3 = ((!(b3-b0))*(p6&&p8));
  assign y4 = (~{{(!(p2?p3:p8))},{4{{p6,p10,p12}}}});
  assign y5 = (3'd7);
  assign y6 = (^(p6+p17));
  assign y7 = (5'd13);
  assign y8 = {(4'd9)};
  assign y9 = $signed(p10);
  assign y10 = (p16<<p6);
  assign y11 = ((((5'd2 * p8)>>(a1===b0))<({a4,b2}==={b1,a4,b1}))+(({p5}^{p15})>=({b0,b1,a4}!=={a2})));
  assign y12 = (a4!==a2);
  assign y13 = ((b1&a0)!==(6'd2 * b1));
  assign y14 = $signed((!((5'd18))));
  assign y15 = (~(~(+(3'sd3))));
  assign y16 = (($signed(b4)?(3'd6):(a2^a3))?$signed(((2'sd1)>>>(a2?p3:a1))):(3'sd1));
  assign y17 = ({4{p1}}>{3{p13}});
endmodule
