module expression_00195(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((&((-3'sd0)<<<(5'sd14)))||(-(3'd4)))^~({(2'd3),(4'd1),(5'd13)}&&((4'sd3)>=(-5'sd6))));
  localparam [4:0] p1 = {4{{4{(5'd25)}}}};
  localparam [5:0] p2 = ({2{{3{(-2'sd1)}}}}<=(~&(((-4'sd7)>=(-5'sd1))&&((2'd2)?(5'sd7):(5'd4)))));
  localparam signed [3:0] p3 = {((2'd0)>>>{3{(-3'sd2)}}),((-(-2'sd1))!=={(4'sd2),(3'd4),(4'd9)})};
  localparam signed [4:0] p4 = ((4'd13)/(4'd1));
  localparam signed [5:0] p5 = ({(+(5'sd10)),((5'sd13)>=(4'd3))}<<<((&(3'd0))+((3'd7)>(-5'sd0))));
  localparam [3:0] p6 = (((3'd5)^(4'd0))?{1{(-4'sd5)}}:{2{(-3'sd1)}});
  localparam [4:0] p7 = ((((5'sd15)&(-2'sd1))>{4{(3'sd3)}})^(((-3'sd3)>=(2'd0))&((4'sd6)<=(-3'sd0))));
  localparam [5:0] p8 = (4'sd6);
  localparam signed [3:0] p9 = ((((-2'sd0)?(5'd5):(5'sd11))>{2{(3'd1)}})==={2{{4{(-3'sd0)}}}});
  localparam signed [4:0] p10 = {(2'd1),{{(2'd3)}},{(+(2'sd0))}};
  localparam signed [5:0] p11 = {{(5'sd6),(4'sd7)},((5'd23)?(4'd11):(2'sd1)),{((4'd4)?(3'd6):(2'd3))}};
  localparam [3:0] p12 = (|(!(5'sd0)));
  localparam [4:0] p13 = ((-3'sd2)>>>(5'sd11));
  localparam [5:0] p14 = (|(+(~^(((-(5'd18))+(!(5'sd0)))!=((^(4'd1))+((3'd3)^~(4'sd2)))))));
  localparam signed [3:0] p15 = (~&(~&(~|{(~|((5'd10)==(5'sd15))),({(4'd2),(-3'sd2)}>>>(&(2'd2))),(!(|(~&(4'd15))))})));
  localparam signed [4:0] p16 = {(((2'd3)?(-4'sd5):(-3'sd1))==((5'd14)^~(-3'sd2))),(((4'd9)&(-5'sd0))?((-3'sd1)?(-2'sd0):(2'sd0)):(+(3'd1))),(6'd2 * ((4'd4)&(4'd3)))};
  localparam signed [5:0] p17 = (5'd2 * ((3'd6)===(4'd13)));

  assign y0 = (((&p11)?(a0?b5:p14):(b2?p14:p4))?((&p14)?(-a4):(~^p9)):((~a5)?(p7?p14:p8):(~a1)));
  assign y1 = ((~(&((+(b0==a2))|(a2+b4))))<<(((~^a0))%b2));
  assign y2 = {(a4&a0),(b1?b1:a5),(p9?p10:p4)};
  assign y3 = ((((b1!==b2)===(a1||b0))<<((b3|p14)>=(b4^~b0)))<<<(((b2<<<b0)==(a5>a3))|{(a3>>>b0),(a0|b4)}));
  assign y4 = (3'sd0);
  assign y5 = {{1{$signed((5'sd0))}},{{1{((~&p1)<<(~|p6))}}}};
  assign y6 = ((~&(p3?a2:p3))||(&(p3-p15)));
  assign y7 = (~^$unsigned((^({{{(2'd1),(+p8),(3'd6)},((+(p14?p9:a3))>(^(a3?a3:p17)))}}))));
  assign y8 = ((|((&(~|a3))>>(~|(2'd0))))<<<(4'd0));
  assign y9 = {{(a4>>b3),(b2|a2),({b4,b2,a2})}};
  assign y10 = {(+((&((|(a3>=b2))|(|{p10})))<$signed((-((~|b0)&&(^b5))))))};
  assign y11 = (~(6'd2 * (a1===b1)));
  assign y12 = (({4{p3}}&&{2{a4}})||({1{({4{p12}}>$signed(a2))}}));
  assign y13 = ({((p10<p2)>>(-(p0&&p16)))}>>>((p9<<<p9)?(p13<=p10):(p13?a3:p11)));
  assign y14 = (2'd0);
  assign y15 = (p4<<p12);
  assign y16 = {2{b1}};
  assign y17 = {1{(~&(|$unsigned((~&{2{{2{p2}}}}))))}};
endmodule
