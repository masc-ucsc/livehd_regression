module expression_00009(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{((2'sd1)!=(-3'sd0))}};
  localparam [4:0] p1 = (3'd2);
  localparam [5:0] p2 = {(5'sd5),(4'd11)};
  localparam signed [3:0] p3 = (&(3'd2));
  localparam signed [4:0] p4 = ((-3'sd1)/(-3'sd2));
  localparam signed [5:0] p5 = (5'd15);
  localparam [3:0] p6 = ({3{(4'd5)}}||{1{((4'd12)<=(5'd1))}});
  localparam [4:0] p7 = (2'sd0);
  localparam [5:0] p8 = ((((-2'sd0)?(-3'sd0):(2'd2))<=((-5'sd9)<<(4'd3)))?(((3'd4)?(4'd4):(3'd5))?((-3'sd2)?(-2'sd0):(2'd0)):((-2'sd0)%(-2'sd0))):(((3'd1)?(3'd3):(5'd4))<<((-4'sd0)&(2'd3))));
  localparam signed [3:0] p9 = (~|{(^(3'd3)),((4'd10)?(-5'sd2):(5'd16))});
  localparam signed [4:0] p10 = (5'sd3);
  localparam signed [5:0] p11 = (((-((5'd18)!==(-4'sd0)))^(+(~|(-3'sd2))))>({3{(3'd2)}}|((5'd17)<<<(-5'sd4))));
  localparam [3:0] p12 = {(!{{(3'd0),(3'd3)},(~&(3'd5)),(-(-3'sd1))}),(+(~^(&(+(+(~^(2'sd0)))))))};
  localparam [4:0] p13 = (4'd11);
  localparam [5:0] p14 = (^(^(~(-3'sd3))));
  localparam signed [3:0] p15 = (|(3'sd3));
  localparam signed [4:0] p16 = (({4{(3'd4)}}==((5'sd8)&(-2'sd1)))>>(5'sd13));
  localparam signed [5:0] p17 = (((3'sd0)&(2'd1))<<(-(-4'sd7)));

  assign y0 = (((2'sd1)!==((a5>>b0)|(a1<=a3)))>(({1{a2}}>>{3{a2}})|((3'sd0)<{1{a4}})));
  assign y1 = (~|(((a3&b2)===(~^b1))>(+{1{(a5|a2)}})));
  assign y2 = ((p3^~p17)&&(|(p8&&b2)));
  assign y3 = {{((a0|b4)===(b3|b4)),({p10,b5}|(p10<p7))}};
  assign y4 = {($unsigned({a2,b2,b5})^~{(a3^b1),(5'd2 * a0)})};
  assign y5 = {a3,p4};
  assign y6 = ($signed(((b1?a2:a4)?(b1?b3:a3):$signed(a5)))!==((|{2{a2}})^~(&(b5?b1:b1))));
  assign y7 = (((~&{p10,a4})));
  assign y8 = (+(~|(|((|(a4&p15))?(b4===a2):(+(b5+b4))))));
  assign y9 = ((4'd2 * (b0^~b0))<=(6'd2 * (b1*a1)));
  assign y10 = $signed({2{p2}});
  assign y11 = (+(~(|(4'd2 * {1{(b0&&p0)}}))));
  assign y12 = (+(~|(({4{a3}}&{1{(b1>>a3)}})<((a0^a1)!=(~|(b4>>>b4))))));
  assign y13 = (((6'd2 * p12)?(a3|p3):(2'd1))>>>(3'd6));
  assign y14 = (~|(~^(-5'sd13)));
  assign y15 = (-(((!(~p15))?((~a5)):(p6?p1:p15))));
  assign y16 = (+(((&p11)?(|p10):(~^p10))?((&p4)?(p17?p1:p1):(p4?p13:p9)):(-((^(a1?b4:a5))===(~&(~|b0))))));
  assign y17 = ({1{((b0>>a1)&&{1{p6}})}}==((~b1)&&{4{a1}}));
endmodule
