module expression_00534(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{{(^((5'd1)>>(5'sd2)))}});
  localparam [4:0] p1 = (5'd27);
  localparam [5:0] p2 = (5'sd11);
  localparam signed [3:0] p3 = {((~^(3'd3))>((3'sd1)+(2'sd0))),{{(-2'sd1),(2'd1),(5'd13)}}};
  localparam signed [4:0] p4 = {2{(|{3{((2'd2)^~(5'd5))}})}};
  localparam signed [5:0] p5 = {3{((-4'sd0)>>>(2'sd1))}};
  localparam [3:0] p6 = {4{{2{(-5'sd14)}}}};
  localparam [4:0] p7 = (2'd0);
  localparam [5:0] p8 = (^(-{((2'sd0)>>(3'sd3)),((2'sd0)!==(3'd6))}));
  localparam signed [3:0] p9 = (&(((5'sd12)^(2'sd1))?(~(-4'sd3)):((4'sd1)?(5'd16):(2'd1))));
  localparam signed [4:0] p10 = ({((2'd0)>>>(2'd1)),((3'd2)>(3'sd2)),((4'sd4)^~(2'd1))}>>>(((5'd16)>>(-2'sd0))==((5'sd10)===(-4'sd5))));
  localparam signed [5:0] p11 = (((4'sd7)===((5'd26)^~(-3'sd2)))===(-2'sd0));
  localparam [3:0] p12 = (((5'd13)?(4'd9):(3'd0))?((-2'sd0)?(-2'sd0):(-4'sd7)):(((-2'sd1)?(-3'sd1):(3'sd3))>=((5'sd7)!=(4'd12))));
  localparam [4:0] p13 = {3{{(2'd1)}}};
  localparam [5:0] p14 = ({(+(3'd4)),((2'd0)^(3'd0))}!==(+(3'd7)));
  localparam signed [3:0] p15 = (4'sd3);
  localparam signed [4:0] p16 = (((2'd0)^~(2'sd1))-((-2'sd0)>=(3'd2)));
  localparam signed [5:0] p17 = ((-{((3'd5)^~(3'd6)),{((3'sd2)&&(3'sd3))}})^~(~^((!((2'sd0)>>>(4'd15)))|(5'd5))));

  assign y0 = ((a3?b1:a5)>>>(~b2));
  assign y1 = (2'sd0);
  assign y2 = (!(-3'sd2));
  assign y3 = (((a3<p13)^(b3?p12:p16))>((p12>>>a4)?(b3?a3:b4):(a2?p8:a4)));
  assign y4 = ((-(p15!=b1))<<{b1,b2});
  assign y5 = (($signed((b2!=b2))&&((b2|b0)))!==((6'd2 * a0)!==(b3?a3:a2)));
  assign y6 = {3{{(3'd3)}}};
  assign y7 = ((~|{4{{p3}}})^~(((^b1)<<<(p3==a5))-{(5'd16),(b2|p7),{p7,p10}}));
  assign y8 = (~(&({(2'd2),(a0|b2)}-({a3,a2,a5}^~(~^b2)))));
  assign y9 = $unsigned({1{$unsigned((((b2>>b0)^(b5<<b0))))}});
  assign y10 = (p12?a3:a0);
  assign y11 = ((a5/b2)==(a3<<a3));
  assign y12 = (((4'd11)>(4'd1))===({(2'd3)}<(5'd2 * b0)));
  assign y13 = ((a0&p4)>=(p16^~p16));
  assign y14 = {1{(((p16&p5)?(b5^p13):{3{p7}})>>>{2{(b1<<p17)}})}};
  assign y15 = ({p16,p7}?$unsigned(a2):(~&p17));
  assign y16 = ((2'd2)<(p9<=p10));
  assign y17 = {4{(~&b5)}};
endmodule
