module expression_00975(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(-((((5'd8)^(5'd19))^~((-5'sd10)&&(-3'sd0)))&(|((2'sd0)+(2'sd0))))));
  localparam [4:0] p1 = (((4'sd1)^~(3'd2))?((-2'sd0)>(3'd6)):(3'd2));
  localparam [5:0] p2 = {((4'd12)&&(2'd0))};
  localparam signed [3:0] p3 = (((+((3'd3)>=(5'sd14)))<={1{((4'sd7)?(-4'sd6):(3'd5))}})!==(~(((5'd17)?(5'sd7):(5'd18))?(~|(3'd5)):((2'd2)?(-2'sd0):(3'sd0)))));
  localparam signed [4:0] p4 = (((5'd2 * (5'd8))|((4'd11)!=(-3'sd3)))<{4{(3'sd0)}});
  localparam signed [5:0] p5 = ((5'd6)?{(5'sd1),(5'sd9),(-5'sd13)}:(5'd2 * (4'd11)));
  localparam [3:0] p6 = (~|((2'd1)?(3'd0):(4'd10)));
  localparam [4:0] p7 = (^(+(~^(((4'sd1)?(4'd14):(5'd16))%(-3'sd3)))));
  localparam [5:0] p8 = {1{(3'd5)}};
  localparam signed [3:0] p9 = (^(3'd3));
  localparam signed [4:0] p10 = (3'sd0);
  localparam signed [5:0] p11 = (3'd2);
  localparam [3:0] p12 = (((~(-4'sd4))>>{2{(2'd0)}})?(~|((2'sd0)?(5'sd2):(5'sd11))):(((5'd25)+(5'sd2))?(!(-2'sd0)):((4'sd0)?(-4'sd3):(2'd3))));
  localparam [4:0] p13 = ((|(|(3'd4)))|((-5'sd2)||(4'sd1)));
  localparam [5:0] p14 = ((^(-(4'd0)))?(~&(~&(4'sd5))):((3'd3)?(-4'sd0):(4'd5)));
  localparam signed [3:0] p15 = {{(^(~&(&(3'd7))))}};
  localparam signed [4:0] p16 = ((2'd2)?(2'sd1):(3'd7));
  localparam signed [5:0] p17 = {(-4'sd5),(((2'd1)+(3'd5))<<(3'd0)),(+(~&(-4'sd2)))};

  assign y0 = (~(~^((^(~p16))^(~|(-p10)))));
  assign y1 = {2{{2{a4}}}};
  assign y2 = (~$signed({4{(|a1)}}));
  assign y3 = (-4'sd4);
  assign y4 = ({{((a1^~p17)||(p5==p4))}}^($unsigned((+p6))!=(~^{p8,a1})));
  assign y5 = (~{{(((-(p2))<<$signed((p14&p11)))||{$signed(p16),(^p15),{b0}})}});
  assign y6 = ({((b3<a3)>={b0,b5,p10}),({4{p10}}?(-2'sd1):(5'd2 * b1))}||{3{(a5?p6:a4)}});
  assign y7 = (!(!(&(~((p10^~b1)>>(+b1))))));
  assign y8 = ((^(4'd12))===(4'd0));
  assign y9 = (!(-(~&(~^(+(&(~(~(|(|(+(~|b1))))))))))));
  assign y10 = ({p9,b3,p9}==($unsigned(p15)<<$signed(b5)));
  assign y11 = ((3'd4)>{1{(b1<=p2)}});
  assign y12 = {{a1},{2{b2}}};
  assign y13 = $unsigned(((-3'sd2)>>>(-3'sd1)));
  assign y14 = $signed(((~^$unsigned((!(|(~&(|p4))))))<$signed((!((~b5)||(!p3))))));
  assign y15 = $unsigned((3'sd3));
  assign y16 = (($signed(a2)!==(b3<b4))>=(5'd2 * $unsigned(b4)));
  assign y17 = ({3{(^{2{p8}})}});
endmodule
