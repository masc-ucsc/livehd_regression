module expression_00287(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({2{(~|(3'd6))}}!=({4{(2'd0)}}===(4'd3)));
  localparam [4:0] p1 = ((-2'sd0)?(2'd1):(5'd27));
  localparam [5:0] p2 = (-(~^(~&(~&(|(~|(3'd1)))))));
  localparam signed [3:0] p3 = (~^{1{(4'sd0)}});
  localparam signed [4:0] p4 = (~(|(-2'sd1)));
  localparam signed [5:0] p5 = (-5'sd0);
  localparam [3:0] p6 = {4{(3'd4)}};
  localparam [4:0] p7 = (((-2'sd0)?(5'd27):(-2'sd1))||((3'd5)+(-4'sd5)));
  localparam [5:0] p8 = ((-2'sd1)?(2'sd0):(3'd4));
  localparam signed [3:0] p9 = (((-5'sd0)?(-3'sd0):(2'd2))?((-5'sd15)?(5'd10):(4'd1)):((5'sd7)>>(2'd0)));
  localparam signed [4:0] p10 = (((-3'sd3)&&(-2'sd0))||((5'sd11)&&(4'sd0)));
  localparam signed [5:0] p11 = ((3'd1)?(~((5'sd15)?(-3'sd0):(-4'sd5))):(((3'd5)?(5'd21):(5'sd7))>>((3'sd3)^(4'sd4))));
  localparam [3:0] p12 = (4'sd5);
  localparam [4:0] p13 = ((((-4'sd1)&(5'sd12))?((-5'sd2)|(4'sd1)):((-5'sd12)<(2'sd0)))==(((3'sd0)&&(-5'sd2))-(4'd2 * (3'd2))));
  localparam [5:0] p14 = (&((^(-5'sd6))==(((4'd8)<=(5'sd2))+((5'sd0)<<<(3'd7)))));
  localparam signed [3:0] p15 = ((&(-5'sd1))?(2'd1):{(3'd3),(4'sd1),(-3'sd3)});
  localparam signed [4:0] p16 = ({((4'd12)?(4'd0):(2'sd1))}?{{(2'd0),(4'd13),(2'sd0)}}:(((3'd7)?(2'sd0):(5'd10))?{(-4'sd7),(3'd0)}:{(5'd27)}));
  localparam signed [5:0] p17 = (3'sd0);

  assign y0 = $unsigned((((3'd6))^~(a0||p9)));
  assign y1 = {2{((+b2)<<{b3})}};
  assign y2 = (~&(5'd14));
  assign y3 = ({3{(p14!=a1)}}?{2{(p6>=p1)}}:$unsigned(((a1?p13:p8))));
  assign y4 = ($signed((a4<b3))?(b2?p17:p1):(4'd6));
  assign y5 = (~(&({(~^(a4+a2)),(|(-a5)),(b4==b3)}-(!(^(+(+(|{(&(a2>=a2))}))))))));
  assign y6 = (p2?p16:a1);
  assign y7 = ({3{{2{p17}}}}>(|{3{p5}}));
  assign y8 = ((((b5?a3:b0)!==(a3?a5:a4))<<<(|(b1||b2)))<=({(a0?p1:a2)}-{{a5,b3,b0}}));
  assign y9 = {3{({(|(a5))})}};
  assign y10 = (4'd11);
  assign y11 = (+(((p16^~a4)>(~(a2?p13:b3)))!=((p3+p2)?(!b0):(p4>>>a3))));
  assign y12 = $signed((({(a1),(~&a0)}!==({b4,b5,a4}))<<<{{4{b1}},$signed((|p17)),((&b3))}));
  assign y13 = {{3{a2}},{4{b1}}};
  assign y14 = $signed(({{a1,b0,p4},$signed({a3,b0,p14})}^~({3{(b4>>>a0)}})));
  assign y15 = {2{(-4'sd3)}};
  assign y16 = {({(a0^~b1),(a1===b4),{a2}}<<<{{p3,a0,b4},{b5}})};
  assign y17 = (^(-(5'd24)));
endmodule
