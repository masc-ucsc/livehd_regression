module expression_00416(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd2)&(5'sd8));
  localparam [4:0] p1 = ((&(((2'd3)+(2'd2))>((5'd11)!=(2'sd1))))<<((((-3'sd3)==(-3'sd2))!==((4'd9)&&(3'd6)))&&(~|(+(~&(-2'sd0))))));
  localparam [5:0] p2 = {{{2{{((-5'sd5)||(5'sd14))}}},{{1{(4'd5)}},{(3'd7),(-2'sd0),(2'd1)},{1{(3'd5)}}}}};
  localparam signed [3:0] p3 = {(2'sd1),(2'd0),(3'sd0)};
  localparam signed [4:0] p4 = ((((2'd0)%(5'sd10))<<<((4'sd2)?(-2'sd1):(3'd0)))<=((4'd6)?(-2'sd0):(-5'sd6)));
  localparam signed [5:0] p5 = (((+(4'd2))<=((-2'sd1)&(-4'sd0)))^~((~^(5'd9))|(~(-2'sd0))));
  localparam [3:0] p6 = (~(2'd3));
  localparam [4:0] p7 = (3'd6);
  localparam [5:0] p8 = {{1{{4{(4'd15)}}}},((4'd2 * (2'd1))?((5'd29)<(3'd2)):((-5'sd10)-(2'd1)))};
  localparam signed [3:0] p9 = {{(-5'sd8)}};
  localparam signed [4:0] p10 = (~^(5'd28));
  localparam signed [5:0] p11 = (({3{(3'd5)}}<<{2{(4'sd1)}})!=({(4'd9),(-3'sd2)}^(|(2'sd0))));
  localparam [3:0] p12 = ((((5'sd7)?(-4'sd1):(-4'sd0))&(~(5'sd14)))!=(((3'd3)?(5'd10):(3'd2))^~((-2'sd0)|(-4'sd7))));
  localparam [4:0] p13 = {(2'd3)};
  localparam [5:0] p14 = {(^(-2'sd0)),(4'd8)};
  localparam signed [3:0] p15 = (+{(3'd1),(4'sd5)});
  localparam signed [4:0] p16 = (((4'sd3)+(-5'sd2))+((-3'sd3)>=(-2'sd0)));
  localparam signed [5:0] p17 = {3{((5'sd13)>>>(4'd14))}};

  assign y0 = ((|$unsigned(($unsigned((a1+a3))>>{(b2||b5)}))));
  assign y1 = $unsigned(((b3?b4:p12)!=(4'd8)));
  assign y2 = (((b2<<p1)>>(p1))?((!a1)?(~|p0):(b0)):(+$signed((-$unsigned(a4)))));
  assign y3 = {1{(~^{4{p8}})}};
  assign y4 = (3'd5);
  assign y5 = (~|(3'd2));
  assign y6 = {1{($unsigned($signed({1{{({{{3{a1}},(~^(&a1)),$signed((+a5))}})}}})))}};
  assign y7 = ((p11/p17)%b3);
  assign y8 = (-4'sd1);
  assign y9 = (-$unsigned({3{({2{$signed(b5)}})}}));
  assign y10 = $signed({2{(!(&{a2,p8,b1}))}});
  assign y11 = (({3{(a4!=p17)}}<<<$signed((~&((b4>>>a2)===$unsigned(b2))))));
  assign y12 = {1{$unsigned({4{(b1)}})}};
  assign y13 = {3{(2'sd1)}};
  assign y14 = (a1^~p7);
  assign y15 = (~&{1{(({1{a2}}^(b4==a5))^((p0<p17)!=(-a5)))}});
  assign y16 = (a5>>a5);
  assign y17 = (-(4'd2 * {2{p14}}));
endmodule
