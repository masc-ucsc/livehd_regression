module expression_00646(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd3)?(4'sd4):(4'd7))?((2'sd1)|(2'sd0)):((-4'sd7)==(5'd30)));
  localparam [4:0] p1 = ((-4'sd2)>=(4'd15));
  localparam [5:0] p2 = ((4'd9)<((4'd0)<<(5'd4)));
  localparam signed [3:0] p3 = ({((5'sd10)&(-4'sd0))}-{1{((4'sd1)!==(4'd4))}});
  localparam signed [4:0] p4 = (~&({(-2'sd0),((3'd6)+(3'sd0)),((2'd3)-(2'sd0))}!==(5'sd3)));
  localparam signed [5:0] p5 = ((((2'd1)<((3'd2)||(3'sd2)))<=(5'sd14))<((|((2'sd1)&&(3'd4)))&(((2'd3)%(-4'sd3))>>(3'sd0))));
  localparam [3:0] p6 = {2{{2{(6'd2 * (|(2'd3)))}}}};
  localparam [4:0] p7 = ((|(((3'd1)>(3'd5))>((2'd2)<<<(4'sd0))))&&(5'd2 * ((2'd1)>>>(5'd29))));
  localparam [5:0] p8 = {{2{((+(2'sd0))<<{2{(4'd12)}})}}};
  localparam signed [3:0] p9 = ((4'd2)?(2'd1):(-3'sd1));
  localparam signed [4:0] p10 = ({1{(&(3'sd3))}}^{3{(5'd17)}});
  localparam signed [5:0] p11 = (-4'sd1);
  localparam [3:0] p12 = ((6'd2 * ((3'd7)<(2'd3)))=={{(-4'sd2),(4'sd0),(5'd8)},(+{(4'd15),(5'd28),(2'd1)})});
  localparam [4:0] p13 = {(3'd6),(-4'sd1)};
  localparam [5:0] p14 = (((4'd10)?(4'sd0):(4'd4))?((4'd15)?(3'd5):(4'd4)):((-4'sd6)?(5'd15):(3'd7)));
  localparam signed [3:0] p15 = {(+(-(!{1{((3'd7)>(2'sd1))}}))),{3{{(-2'sd0),(5'd29)}}}};
  localparam signed [4:0] p16 = (&(((-3'sd0)?(4'd12):(3'sd2))>(!(|(3'sd0)))));
  localparam signed [5:0] p17 = {({3{(3'sd2)}}>>(+((3'sd1)>>>(4'sd1)))),(~^{3{(+(2'sd1))}})};

  assign y0 = ({2{($unsigned(a1)-(b0<b1))}}|{(!(b5)),$signed((b4)),{3{a1}}});
  assign y1 = {4{(2'd0)}};
  assign y2 = (&$signed({(+(($unsigned(b4)))),((~|(p3?a0:a5))),((p0?a2:p4)>>>(-a1))}));
  assign y3 = (3'd1);
  assign y4 = {1{((&(~|(-(p2?p15:b1))))?(^(~{3{p14}})):(~&(|(~^(&{1{p11}})))))}};
  assign y5 = ((+(+((p13^p15)?(a1^b4):(p7+b3))))+(($signed(a1)!=(p6?p0:p16))&((p16-a4)!=(b0>>>b2))));
  assign y6 = $signed(((~(~|(+(~(p0^~b1)))))<<<(-4'sd5)));
  assign y7 = $signed({{{b2},(p9),(p2!=p13)}});
  assign y8 = {4{b2}};
  assign y9 = (p3?p16:p3);
  assign y10 = $signed((2'd3));
  assign y11 = (~|{$unsigned(((6'd2 * p12)-(5'd2 * b0))),$unsigned(((p5||a5)==$signed(p4)))});
  assign y12 = (b1?a4:p17);
  assign y13 = {((p7<<<p7)&{p10}),(-2'sd0)};
  assign y14 = (+{{(p5),{p2,p12},(p17)},{(p2>p9),(~|$signed(p3))}});
  assign y15 = (~&(5'd22));
  assign y16 = ((~|b5)<(b5!==a3));
  assign y17 = (p10?p11:p9);
endmodule
