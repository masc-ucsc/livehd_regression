module expression_00743(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((3'sd1)?(+{4{(4'd2)}}):(+((4'sd7)?(5'd20):(-4'sd0))))};
  localparam [4:0] p1 = ((((2'd1)==(3'sd3))>{3{(2'sd0)}})===({2{(-2'sd0)}}>>((4'd12)!==(3'sd1))));
  localparam [5:0] p2 = ((((4'd15)>(-4'sd7))===((-3'sd1)?(5'd4):(3'sd2)))?(+(-((2'sd1)?(5'd4):(3'd1)))):(((-3'sd3)!==(-3'sd1))==((2'd1)?(5'sd3):(4'd0))));
  localparam signed [3:0] p3 = ((((-2'sd1)^~(-2'sd1))?((3'd2)>>(-3'sd3)):((3'd0)<=(3'd1)))===(((-4'sd6)===(4'd12))+((-2'sd1)+(-3'sd0))));
  localparam signed [4:0] p4 = ((-(|(~|(-2'sd0))))?{(~^(~^(4'd6)))}:((4'sd1)?(-4'sd1):(5'sd12)));
  localparam signed [5:0] p5 = (^{1{(4'sd4)}});
  localparam [3:0] p6 = (&(~|(((~(4'sd5))>>(~^(5'd12)))<=(|(~(+(~&(4'd8))))))));
  localparam [4:0] p7 = (-(3'sd3));
  localparam [5:0] p8 = (((4'sd6)?(5'sd9):(4'd2))===((4'd7)<<(5'd29)));
  localparam signed [3:0] p9 = (((4'd4)?(-3'sd3):(2'd2))?((-3'sd1)!==(3'd7)):{(-(3'sd0))});
  localparam signed [4:0] p10 = (((+((-5'sd3)!==(3'sd2)))!==((5'd31)&&(2'd1)))>=(((2'd0)?(2'd0):(3'sd0))?(+(4'sd0)):(~(5'd23))));
  localparam signed [5:0] p11 = (|(^(~&((3'sd3)==(^((3'd1)/(-2'sd1)))))));
  localparam [3:0] p12 = ((((2'd2)===(-5'sd1))/(5'sd15))^(4'd3));
  localparam [4:0] p13 = ((+(-(^((4'd1)?(-2'sd1):(-5'sd6)))))?(((3'd1)|(3'd3))-((5'd22)||(3'd6))):((|(4'd7))>((3'd0)?(-5'sd3):(-4'sd7))));
  localparam [5:0] p14 = ((((4'd9)||(5'd29))||((3'sd0)>>>(5'd4)))+(((3'sd2)-(3'd1))>>>(!(2'sd0))));
  localparam signed [3:0] p15 = ((4'd12)?(2'd0):(-5'sd2));
  localparam signed [4:0] p16 = ((4'd3)>>>(3'd4));
  localparam signed [5:0] p17 = ({3{((-5'sd5)?(5'd10):(2'd3))}}&(6'd2 * ((3'd3)>>>(5'd23))));

  assign y0 = {1{(4'd2 * (^(6'd2 * p8)))}};
  assign y1 = {3{p2}};
  assign y2 = (-5'sd6);
  assign y3 = ((~|(a1&&a1))<(~(p3<<<b5)));
  assign y4 = ($signed((|(($signed((|($unsigned(a2)&(-2'sd1)))))^~({4{b3}}<(a5|b0))))));
  assign y5 = (|(a4>=a4));
  assign y6 = ({2{p17}}!=(~|{4{b3}}));
  assign y7 = (&(b4>>>a0));
  assign y8 = (&(&$unsigned(p13)));
  assign y9 = ((2'sd0)?((+a3)?(b1?p7:b5):(-3'sd0)):((&a1)?(a1):(~&p6)));
  assign y10 = (-4'sd6);
  assign y11 = ({4{p15}}?{p12,a3,p8}:(p4<=a3));
  assign y12 = (b4||a5);
  assign y13 = ((b1/b0)<(|(p13?b4:a5)));
  assign y14 = (($signed($unsigned((b2+b3)))===$signed(({4{b4}}<(-5'sd1))))!==(3'sd2));
  assign y15 = (p15<<<p1);
  assign y16 = {{3{{2{a1}}}},(4'd8)};
  assign y17 = (({3{b4}}&{b0,b1,b5})|(((a1>>>a4)===(b3^~b3))>>((p17|p17)<<<(p2<<b3))));
endmodule
