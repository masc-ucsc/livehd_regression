module expression_00840(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd7)||(3'sd2))<(+(4'd12)));
  localparam [4:0] p1 = (~|(~&{1{(-(~|((-5'sd1)?(-4'sd0):(4'sd4))))}}));
  localparam [5:0] p2 = (((3'd3)?(2'd2):(-4'sd2))?(4'd2 * (+(4'd5))):(-5'sd8));
  localparam signed [3:0] p3 = {{(-4'sd1),(-3'sd1),(-2'sd0)},{(4'd11),(3'sd3),(-4'sd6)},{(4'sd3)}};
  localparam signed [4:0] p4 = (4'd2 * ((2'd2)?(3'd1):(4'd9)));
  localparam signed [5:0] p5 = {(4'sd5)};
  localparam [3:0] p6 = (-4'sd3);
  localparam [4:0] p7 = (+(-2'sd0));
  localparam [5:0] p8 = {(-4'sd3),(2'd0),(5'd26)};
  localparam signed [3:0] p9 = {2{(3'd6)}};
  localparam signed [4:0] p10 = {1{{{3{(2'd2)}},((4'd2)?(4'sd4):(5'd17))}}};
  localparam signed [5:0] p11 = ({((4'd10)-(-5'sd6)),((4'd4)<=(5'sd9))}^(^(((5'd5)^~(3'd2))&{4{(-4'sd6)}})));
  localparam [3:0] p12 = {4{(4'd12)}};
  localparam [4:0] p13 = {4{((3'sd1)===(4'd11))}};
  localparam [5:0] p14 = ((&(-2'sd1))?(~&(5'sd10)):((2'sd1)==(5'd4)));
  localparam signed [3:0] p15 = ((-5'sd12)>>>(3'sd0));
  localparam signed [4:0] p16 = (&({(^(4'd4)),(~&(5'd29))}?{(|{(2'sd1),(-5'sd1)})}:((-4'sd3)?(5'd12):(-3'sd3))));
  localparam signed [5:0] p17 = {(|(5'sd15)),{(5'd3),(3'd4)},(-3'sd1)};

  assign y0 = ((5'd22)?(+(a3?b3:a5)):(-(4'd13)));
  assign y1 = (((4'd4)?(a5-p4):{4{b5}})!=(3'd3));
  assign y2 = (~^(~&(~|(~|(!(&((~(a3||b2))-(!{2{p14}}))))))));
  assign y3 = {4{(a1|p13)}};
  assign y4 = (-4'sd1);
  assign y5 = (~&b0);
  assign y6 = ($unsigned({{b3},{a0,p15}})?$unsigned($unsigned((~|(p13<=p10)))):(3'sd1));
  assign y7 = ((((p13+p0)^~(p9==p17))>((b2!==a2)>(p10>>p14)))!=(((b0||a1)>=(b3>=b3))===((b0+b5)&(b1!==b2))));
  assign y8 = {4{(3'd0)}};
  assign y9 = (2'd2);
  assign y10 = (~|(((!(p16&b2))<<<(2'sd0))!=((~(p16-a0))<{1{{p8,p11}}})));
  assign y11 = ((a5)<(~|p16));
  assign y12 = ((&(~&((~|(p11&p8))<=(-(a1-b0)))))||(~|(~^((p5&&p8)<=(~|(p3<<b1))))));
  assign y13 = (+(4'd1));
  assign y14 = {(4'd4)};
  assign y15 = (6'd2 * (p6&&p2));
  assign y16 = $unsigned((($unsigned(b1)||(p2))>>>((a4)?(b5>=a1):(p13?p4:a3))));
  assign y17 = (5'd14);
endmodule
