module expression_00275(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(4'd10));
  localparam [4:0] p1 = ((-2'sd1)?(4'd6):{2{((-5'sd12)!=(3'sd3))}});
  localparam [5:0] p2 = (-5'sd0);
  localparam signed [3:0] p3 = (~&((+((-4'sd0)%(2'd3)))<(~|(^((2'd0)<=(-2'sd0))))));
  localparam signed [4:0] p4 = (((^(-5'sd5))&&(|(4'd1)))^(6'd2 * ((3'd7)<(2'd0))));
  localparam signed [5:0] p5 = {4{(2'sd0)}};
  localparam [3:0] p6 = (((2'sd1)^~(4'd14))/(5'd30));
  localparam [4:0] p7 = {1{((2'd0)|(5'sd4))}};
  localparam [5:0] p8 = {1{{(4'd10),(5'sd7)}}};
  localparam signed [3:0] p9 = {(({(5'd26),(4'sd7)}+{(4'sd5),(5'd12)})+({(3'd1),(5'd14)}?((2'd2)?(5'd20):(3'd4)):((-5'sd7)<<(-3'sd2))))};
  localparam signed [4:0] p10 = ((3'd7)|(3'sd3));
  localparam signed [5:0] p11 = (((3'd5)<<(4'd0))!=((2'sd0)>>>(3'd3)));
  localparam [3:0] p12 = (~^((|(2'd3))<<<{2{(2'd0)}}));
  localparam [4:0] p13 = ((((4'd1)>>>(4'd7))>=(~&(2'sd0)))||((-(5'd19))<<<((3'd1)>>(4'd12))));
  localparam [5:0] p14 = {(2'sd0)};
  localparam signed [3:0] p15 = ({(5'd29),((3'd1)&(-4'sd6)),((-5'sd13)<<<(2'sd0))}^{2{(2'sd1)}});
  localparam signed [4:0] p16 = {{(((4'd15)|(2'sd1))<((4'd8)<(2'd1)))},(^{{(3'd7),(-2'sd0)},((-2'sd1)?(-3'sd0):(4'd6))}),(+{(~{(-3'sd0)})})};
  localparam signed [5:0] p17 = (|{(5'sd4),(5'sd14)});

  assign y0 = ((^p16)?(3'd5):(-3'sd0));
  assign y1 = (~^(!(5'sd6)));
  assign y2 = (&(+$signed(((((-b2)^~(b5))&&((~&b5)/b1))>>>((!(b5&b1))==$unsigned(((~|a2))))))));
  assign y3 = (4'sd7);
  assign y4 = (-2'sd1);
  assign y5 = ({4{(b4<<<p1)}}<((p14>=b0)<<<(b1!==a2)));
  assign y6 = {2{{2{(4'd7)}}}};
  assign y7 = (&(~$unsigned((b4==a0))));
  assign y8 = (5'd21);
  assign y9 = (6'd2 * {(b2|p7)});
  assign y10 = (((b4<<b4)>>>(~(a2!==b2)))^((4'd2 * (p1|a1))));
  assign y11 = ({1{{3{(b3-a5)}}}}?((a1!=a3)?{2{b1}}:$signed(a4)):({3{a4}}?(a5^b5):(b4)));
  assign y12 = (({4{p7}}?(p2<<<p0):{3{p8}})>>>(5'd5));
  assign y13 = $signed(a4);
  assign y14 = ($unsigned((((a3?a2:a5)^(a1&&a1))))>>{1{((b3)<={4{p8}})}});
  assign y15 = ($signed((~(&(((+b5))?(!(b3?b3:a0)):(|$signed(a4)))))));
  assign y16 = ({1{(|((p12?p14:a3)<=(p16?b4:a5)))}}>>($signed((5'd2 * a1))>>>(~&(&p13))));
  assign y17 = (((b1|b3)?{2{a5}}:(b0-b4))==((b1?p14:b3)-(b1!==b1)));
endmodule
