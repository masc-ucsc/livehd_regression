module expression_00091(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{3{((3'd7)?(4'd0):(5'd15))}}}};
  localparam [4:0] p1 = {(~{(&((3'sd0)>(5'sd1))),(^{2{(-2'sd0)}})})};
  localparam [5:0] p2 = (-(|((-((5'd28)*(4'd11)))!=(~(~&(!(-3'sd2)))))));
  localparam signed [3:0] p3 = ({1{(4'd0)}}>>((4'd13)>=(4'd5)));
  localparam signed [4:0] p4 = (|(5'd2 * (!{1{(5'd26)}})));
  localparam signed [5:0] p5 = ({((-4'sd5)===(-5'sd0))}-((4'd4)>>(-5'sd6)));
  localparam [3:0] p6 = (({2{(2'd3)}}<((2'd1)>(4'd2)))<<(((3'sd2)-(4'sd2))<<<((3'd6)?(-4'sd5):(5'd1))));
  localparam [4:0] p7 = (2'd0);
  localparam [5:0] p8 = (({(-2'sd0),(5'sd3)}<=((-4'sd5)&&(3'd6)))-({4{(3'sd1)}}<((4'd1)<(4'd15))));
  localparam signed [3:0] p9 = ((-((3'd6)?(4'd13):(4'd0)))?((2'd1)!==(2'sd1)):((-2'sd0)-(4'd13)));
  localparam signed [4:0] p10 = (((3'sd0)>>>(-4'sd4))?((2'd0)!=(-4'sd4)):(~|(5'd2 * (4'd13))));
  localparam signed [5:0] p11 = (~^(((+(-5'sd4))<{(4'd3)})===(~&(-((2'd1)|(2'sd1))))));
  localparam [3:0] p12 = (2'sd1);
  localparam [4:0] p13 = {{((-4'sd5)?(2'sd0):(-3'sd1))},((-5'sd14)?(4'd5):(2'sd1)),((-3'sd3)<<(3'sd1))};
  localparam [5:0] p14 = ((4'd2 * (5'd17))>>>((4'd10)<<(-3'sd2)));
  localparam signed [3:0] p15 = (|(+(((5'd28)?(5'd13):(-2'sd0))?(&((3'd6)<(3'd0))):((4'sd6)?(-2'sd1):(-3'sd3)))));
  localparam signed [4:0] p16 = (+((~((5'd9)?(2'd3):(-3'sd2)))?(((-2'sd1)!==(-2'sd0))<<((-4'sd0)>=(-5'sd1))):(((2'd2)?(4'd8):(5'sd8))?((-5'sd11)/(2'd1)):(-3'sd1))));
  localparam signed [5:0] p17 = ((((3'sd0)==(4'd4))>=((3'd1)&(5'd10)))-(((3'd2)!==(-3'sd1))<((-2'sd1)%(3'sd1))));

  assign y0 = ({b0}<=(p0||p7));
  assign y1 = ((&p12)&&(|b5));
  assign y2 = (|(((6'd2 * b0)!==(a4<=b1))>>((&p13)<(p4>>p6))));
  assign y3 = (5'd2);
  assign y4 = {(^(^(-3'sd1)))};
  assign y5 = ({1{b5}}<<<{4{b4}});
  assign y6 = (&((p12?p3:p16)));
  assign y7 = (!($signed((((^a0)?(b1%p16):(a4!=a2))?(~&(^(b0&b1))):((b1?a5:a5)!=(~|a1))))));
  assign y8 = {3{{4{a0}}}};
  assign y9 = (~&(~^(-2'sd0)));
  assign y10 = (!{(-(-(~^{(+{p5,b5}),(!(+b5))}))),{{2{{3{a1}}}},{1{{1{{(~&b1)}}}}}}});
  assign y11 = ((b5||p9)?(~(&p16)):(a2===b5));
  assign y12 = ((p4?b0:a1)?{1{b3}}:(a3));
  assign y13 = ((~^(~^($signed((p6^p15))!=(!$unsigned(p14)))))>>((((~|p12)>>(^p6))|((p4*p5)+(-p9)))));
  assign y14 = (2'sd0);
  assign y15 = {(p16<<p8),(b0^~p8),$unsigned((p15|p11))};
  assign y16 = ((4'd11)?(~|(b0?p7:a5)):$unsigned((!p12)));
  assign y17 = (^((+(2'd3))<=(+((~&(2'sd0))<<<((-2'sd1)>>>(~p13))))));
endmodule
