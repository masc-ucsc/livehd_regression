module expression_00110(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd3),(5'sd8)};
  localparam [4:0] p1 = ((4'd2 * ((4'd13)?(3'd2):(3'd6)))==(|((&((3'd7)&(5'd29)))&((-2'sd0)&&(3'd0)))));
  localparam [5:0] p2 = ({{(3'd2),(2'd1),(5'sd6)}}^~({(3'd3)}&&(6'd2 * (2'd0))));
  localparam signed [3:0] p3 = (&(+(5'd4)));
  localparam signed [4:0] p4 = (-2'sd0);
  localparam signed [5:0] p5 = (+(~|((4'sd5)!=(3'd4))));
  localparam [3:0] p6 = (~^(!(2'd0)));
  localparam [4:0] p7 = (5'd0);
  localparam [5:0] p8 = (-3'sd2);
  localparam signed [3:0] p9 = (^((2'd1)^(((-2'sd1)||(3'd5))|((3'd2)&&(-3'sd3)))));
  localparam signed [4:0] p10 = {({(5'd7),(4'd2)}?{(4'd2),(5'd11),(-5'sd13)}:((3'd5)<<(-5'sd12)))};
  localparam signed [5:0] p11 = {{4{(-2'sd0)}},{1{{{{(-2'sd1)}}}}},{{3{(2'd3)}},{(5'd29),(5'd8)}}};
  localparam [3:0] p12 = (-3'sd0);
  localparam [4:0] p13 = {3{((2'sd1)?(5'd20):(3'sd3))}};
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = (((-5'sd11)<(-3'sd0))^~{3{(3'sd1)}});
  localparam signed [4:0] p16 = (2'sd1);
  localparam signed [5:0] p17 = (((5'sd1)!=(-3'sd0))<=((2'd1)|(-5'sd7)));

  assign y0 = {{(p8<b3)},(a2&p4),{(4'd9)}};
  assign y1 = ((({b2,p12,p8}?(a3<<a5):(~a1))&&((a5?a3:b1)<<(b4?b0:b0))));
  assign y2 = ((4'sd7)||(p4));
  assign y3 = {2{((a3?b1:p1)?{1{b2}}:{2{p0}})}};
  assign y4 = (((2'sd0)^{2{p5}})-((3'd7)==(!p8)));
  assign y5 = ({2{(a4^~b4)}}?{3{(-4'sd5)}}:{3{(b4?a0:a0)}});
  assign y6 = {((a1===a2)&$signed({3{b3}})),({2{a0}}>>>{3{a3}})};
  assign y7 = ((a2?a5:p1)?{b4,a1,b4}:$unsigned(b0));
  assign y8 = (((p3==p2)<(p8/p4))<=(^(&(~((~a1)<(p11*a4))))));
  assign y9 = (|({b2,a4,a5}<(p8>b0)));
  assign y10 = (^((4'sd3)));
  assign y11 = ((4'd2 * (^(p14||p14)))=={3{(&p9)}});
  assign y12 = ((a5+a3)<<<(b4?a1:p0));
  assign y13 = ((((b5^p5)||$signed(p0))&{2{(a4>>>b1)}})<=(^((p2>=p0)|{a3,b1})));
  assign y14 = (4'd8);
  assign y15 = (&({2{{4{a0}}}}>>({2{{2{p6}}}}>>{3{a1}})));
  assign y16 = (2'd3);
  assign y17 = (((~^(p15-p2))?((p4^~p2)):(+(~^p15)))!=(&(~&(~($signed((a0?b2:a3))===(!(-a2)))))));
endmodule
