module expression_00193(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{{(~(!{{(3'd0),(-4'sd0),(3'd4)},{(5'sd13),(2'sd0)},(^(5'd10))})),{{(4'sd0)},(+(-2'sd1)),{(5'd10)}}}}};
  localparam [4:0] p1 = (-4'sd1);
  localparam [5:0] p2 = (~|(&(5'd18)));
  localparam signed [3:0] p3 = (((5'd5)<<<(5'sd1))!==((5'sd0)+(2'd1)));
  localparam signed [4:0] p4 = ((((5'd13)>>(2'd3))&&((5'd21)<=(5'd30)))<(((3'd7)!==(4'sd2))-((4'd10)-(5'd26))));
  localparam signed [5:0] p5 = ((4'd6)<<(4'd5));
  localparam [3:0] p6 = ((!({2{(3'd2)}}>={3{(3'd5)}}))+(|(((4'sd5)?(-5'sd9):(4'd14))&&((3'd2)?(4'd10):(3'd2)))));
  localparam [4:0] p7 = (&(((2'sd1)|(2'd1))*(-((-2'sd0)==(-2'sd0)))));
  localparam [5:0] p8 = (^(~|(5'sd15)));
  localparam signed [3:0] p9 = (+{(({(-3'sd0),(3'd4),(3'd0)}==(~|(2'd1)))?(((4'sd5)?(5'd30):(3'sd1))!=((5'd30)>>(3'd2))):(((4'd14)?(5'd18):(3'd3))!={(3'sd2),(5'd1)}))});
  localparam signed [4:0] p10 = {(!{(|(~{(!(4'd5))})),(!{((4'sd6)===(-3'sd3)),(~(4'sd2))})})};
  localparam signed [5:0] p11 = {2{({3{(4'd13)}}!={2{(2'd3)}})}};
  localparam [3:0] p12 = (~|{(-2'sd0),(3'd1)});
  localparam [4:0] p13 = (-5'sd13);
  localparam [5:0] p14 = (4'd8);
  localparam signed [3:0] p15 = {1{{3{(~^((3'sd3)>>>(2'd1)))}}}};
  localparam signed [4:0] p16 = (3'd6);
  localparam signed [5:0] p17 = (-5'sd8);

  assign y0 = {1{((-5'sd8)>=$signed($signed((~|(~&$unsigned(p15))))))}};
  assign y1 = (~^(((a3===b3)|(~(b4<<<b3)))!==((a4+b0)*(b2+a4))));
  assign y2 = ((a4&p0)<<{{p17,a2,p6}});
  assign y3 = (((+b2)?(a0<<b3):(a4!=b1))===((a0?b1:b1)?(~&a4):(~a3)));
  assign y4 = (2'd1);
  assign y5 = (!((-4'sd1)));
  assign y6 = (({2{p17}}<=((p11||a5)))^~($unsigned((~&a0))<<<(b3>a3)));
  assign y7 = (~&(!(&$signed(((~&(b2<=p13))?(p11?p17:p6):(~$unsigned(b2)))))));
  assign y8 = (((p5?a5:a3)?(b4%a1):(b5?p10:p0))?((p9>>>p10)?(p0?p0:p4):(b1>=a5)):((p12<<p4)&(3'd3)));
  assign y9 = (~(~^(!(~(5'd18)))));
  assign y10 = (3'd2);
  assign y11 = (4'sd5);
  assign y12 = ((p10>>>p10)?(a2===b3):(p3?a1:b2));
  assign y13 = (({b4,a3}^{b3,a1,b4})>>>({1{a2}}?(b1+b5):(p5<<<b2)));
  assign y14 = $signed((({4{b2}})+{2{(b5!=b3)}}));
  assign y15 = (^$signed((~p2)));
  assign y16 = ((6'd2 * a1)<={2{p10}});
  assign y17 = (~((-((4'd2 * {1{(4'd12)}})>{4{{2{a3}}}}))));
endmodule
