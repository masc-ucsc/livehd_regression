module expression_00164(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'sd8)?(4'd1):(4'd10))<(4'd12));
  localparam [4:0] p1 = ({(5'd9),(3'd7)}&{((5'sd6)|(-3'sd2))});
  localparam [5:0] p2 = (4'sd1);
  localparam signed [3:0] p3 = ({3{(2'sd1)}}+{(2'sd1),(5'd1),(4'd8)});
  localparam signed [4:0] p4 = (2'd0);
  localparam signed [5:0] p5 = (^((((2'd0)||(2'd1))?(5'd6):((5'sd15)&(2'd2)))!=({((4'd10)&&(5'sd13))}<<((4'sd7)+(3'd0)))));
  localparam [3:0] p6 = (4'd2);
  localparam [4:0] p7 = {3{((2'd3)>((-5'sd0)>>>(4'd12)))}};
  localparam [5:0] p8 = ((((3'd7)-(5'd3))>=((3'sd3)+(-4'sd6)))<={{(5'd10),(5'd30),(-2'sd1)}});
  localparam signed [3:0] p9 = ((((-3'sd0)?(-4'sd7):(2'sd1))<{3{(2'd0)}})?(((-2'sd1)+(4'd3))?((5'sd4)?(4'd6):(-5'sd1)):((5'd5)?(3'd3):(-2'sd1))):(((-4'sd5)?(-4'sd0):(-3'sd0))?((-2'sd1)<<(2'sd0)):((3'd7)?(-2'sd0):(-2'sd0))));
  localparam signed [4:0] p10 = ((-3'sd2)&&(((3'sd0)>(3'sd3))>=(|(3'd0))));
  localparam signed [5:0] p11 = ((((2'd2)?(-5'sd11):(2'd0))?((5'd25)?(5'sd2):(3'sd0)):((-4'sd2)?(3'd6):(-4'sd4)))===((((3'sd2)<(3'sd2))>>((2'sd0)?(5'd1):(3'd2)))==(((5'd17)?(3'd6):(3'd6))&((2'sd1)>=(5'sd5)))));
  localparam [3:0] p12 = ((((2'd1)!=(2'd2))<=((5'd18)+(-2'sd0)))&(-(~&(!(4'd12)))));
  localparam [4:0] p13 = (3'd0);
  localparam [5:0] p14 = (((((2'sd1)>(-5'sd10))==((-2'sd0)>=(-2'sd0)))>={(-4'sd2),(4'd2),(5'd5)})>>>(((2'd1)?(4'd14):(4'd1))?{(3'd1),(-2'sd0)}:((5'sd12)<<<(-2'sd1))));
  localparam signed [3:0] p15 = (&(~&(3'sd2)));
  localparam signed [4:0] p16 = (((2'd2)&&(2'sd0))==(4'd2 * (5'd26)));
  localparam signed [5:0] p17 = (((5'd24)%(3'd1))<<((2'd0)*(5'sd4)));

  assign y0 = {(2'sd1)};
  assign y1 = (~&(~$unsigned((-(~&p0)))));
  assign y2 = {3{((b0>=a3)>(4'd2 * p14))}};
  assign y3 = ((&((b3?p2:p9)<(a5==p5)))^((-2'sd0)?(a5!==a0):(p6?p9:p5)));
  assign y4 = ((~&(|((b0||p17)^~(~&a1))))<<<((!{b4,p15,b0})-{1{{3{p1}}}}));
  assign y5 = {(p1?p12:p3),(-5'sd5),(p13?p2:p1)};
  assign y6 = (~{((+p17)&(~|p4))});
  assign y7 = ({4{b1}}?((p16?b3:a1)?(a2|a5):{3{p14}}):{3{(b3<a2)}});
  assign y8 = {1{({3{{2{b2}}}}!=={4{{b3,b5,a4}}})}};
  assign y9 = (b2?b4:a1);
  assign y10 = (p6&&a2);
  assign y11 = (5'd2 * (p14&p13));
  assign y12 = ((-{(2'd0)})>{3{(3'd1)}});
  assign y13 = ((((~(^p14))*(&(a1)))));
  assign y14 = (4'd11);
  assign y15 = (((&p3)?(b1^~p7):(-p15))?({p2}?(2'd0):(-2'sd1)):$signed((-(p12?p1:p11))));
  assign y16 = (((p10?a5:p0)&&(a1^a5))?((4'd11)%a0):(-2'sd1));
  assign y17 = ($signed(p1)>=(p0));
endmodule
