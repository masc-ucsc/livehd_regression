module expression_00793(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((|(-5'sd10))||(~^(^(5'd29))))^~(3'd4));
  localparam [4:0] p1 = (!(-4'sd1));
  localparam [5:0] p2 = (4'sd6);
  localparam signed [3:0] p3 = {4{({2{(2'd2)}}===(2'sd0))}};
  localparam signed [4:0] p4 = {((2'sd0)!=(!(((4'd5)!==(-5'sd15))^~{4{(5'd8)}})))};
  localparam signed [5:0] p5 = (-5'sd14);
  localparam [3:0] p6 = {{(^(4'sd7)),{(2'd2)}},(((5'sd10)===(2'd0))^~((-4'sd7)&(4'd15)))};
  localparam [4:0] p7 = (~(-{3{((3'd5)==(3'd7))}}));
  localparam [5:0] p8 = (&((((3'd7)>>>(2'd0))!==(-{(3'd4)}))>>((-(5'd2 * (4'd4)))!=(6'd2 * (3'd0)))));
  localparam signed [3:0] p9 = (((2'd0)>>>(5'd21))?(|(3'sd1)):(~(4'd8)));
  localparam signed [4:0] p10 = ((~^(-2'sd0))?(!(2'd1)):((3'd2)<<(-4'sd2)));
  localparam signed [5:0] p11 = ((+(-2'sd0))?((4'd2)?(2'sd0):(5'd30)):((-2'sd0)?(4'd14):(-3'sd1)));
  localparam [3:0] p12 = ({{((2'd3)?(5'd27):(3'd2))}}>>>(3'd7));
  localparam [4:0] p13 = (~|{2{(|((4'd11)<<(-5'sd12)))}});
  localparam [5:0] p14 = {((~^(3'd0))^(~&(-3'sd1))),(~|({(5'd20),(3'd4)}-{3{(5'd13)}}))};
  localparam signed [3:0] p15 = ((3'd7)&&(4'd10));
  localparam signed [4:0] p16 = (~|((!(((4'd13)>>(-3'sd1))?(-(-3'sd2)):(^(2'd2))))>>(3'sd2)));
  localparam signed [5:0] p17 = {(((5'd26)&&(3'sd0))===((-2'sd1)!=(-5'sd0))),(((5'd4)^~(4'd8))!=((2'd0)!==(5'd22))),{(2'sd0),(3'd1),(2'sd1)}};

  assign y0 = (4'd1);
  assign y1 = (((6'd2 * a2)=={1{a2}})>>{$signed({4{a2}})});
  assign y2 = ((a3>p4)?(^(b0?p2:p15)):(-5'sd14));
  assign y3 = (b4<b4);
  assign y4 = (~|($unsigned(p16)>>>(a0)));
  assign y5 = (!{1{(5'd23)}});
  assign y6 = ($signed(((b4&&b1)&(~|(a2^~b4))))!==(+((!(b5))^~$unsigned((a0<<<a1)))));
  assign y7 = ((({b3,p5,b5}|{3{p4}})>{{b2,b0,p14}})>>((5'd24)?(p15?b3:p17):(b2-p13)));
  assign y8 = (((p3?p6:b3)?(p0<<<b3):((b1)))||({(p15&p0),{b2,b3},(b1!=a3)}));
  assign y9 = ({3{(a1&b2)}}!==({3{a3}}>>>{1{(b4<=a2)}}));
  assign y10 = (p14<<p1);
  assign y11 = (2'sd1);
  assign y12 = ({(a0>>>b2),(|(b0?a5:a4)),$signed((-a5))}===(~^((-(&b5))>>>(-(b5?b1:b4)))));
  assign y13 = (~((!(-(~|(~{p0,p10}))))+((+p8)?(~|p13):(^p10))));
  assign y14 = ($signed((2'sd0))||(^(~^(~^$unsigned((!(^(p3&p9))))))));
  assign y15 = (3'd7);
  assign y16 = (({p3,b5}>=(p1==b3))+((&{a0})));
  assign y17 = (((~^p13)^~(b2^~b4))^~(3'sd0));
endmodule
