module expression_00247(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {({(5'd6)}!==(4'd10)),{(-3'sd0)}};
  localparam [4:0] p1 = (&((|((3'sd2)==(2'd1)))/(3'sd0)));
  localparam [5:0] p2 = (5'sd13);
  localparam signed [3:0] p3 = (~^(!(-((|(5'd9))>>(5'sd12)))));
  localparam signed [4:0] p4 = (((4'd0)?(3'd7):(2'd0))-{(3'd3),(2'd2)});
  localparam signed [5:0] p5 = ((5'd22)?(-3'sd2):(4'sd5));
  localparam [3:0] p6 = ((|(~((~(2'd3))*(-(2'sd1)))))>(~(~&(&(~|(~^((3'sd3)^~(-5'sd1))))))));
  localparam [4:0] p7 = {(+(((3'd1)>{(-4'sd6),(4'sd6),(3'd7)})>>>{(-2'sd1)}))};
  localparam [5:0] p8 = (4'sd4);
  localparam signed [3:0] p9 = (&(~&(-(~^(+(+(|(~^(+(~|(~&(3'd0))))))))))));
  localparam signed [4:0] p10 = (((2'd1)?((3'sd3)?(-4'sd7):(5'd30)):((4'd9)?(4'sd2):(2'sd1)))===(((-4'sd7)<<(5'd16))?((4'd12)&&(-3'sd0)):((-5'sd7)&(5'd23))));
  localparam signed [5:0] p11 = (5'd2 * (~^((4'd9)>>>(5'd10))));
  localparam [3:0] p12 = (((5'sd11)?(3'sd2):(5'sd14))?((4'd0)?(5'd21):(-4'sd5)):(~|(2'd0)));
  localparam [4:0] p13 = (!(~^{(2'd2),(~(+(~&(~&(-5'sd13)))))}));
  localparam [5:0] p14 = (({3{(2'd3)}}?((4'sd3)?(2'd0):(5'd2)):((-2'sd1)?(2'sd0):(5'd20)))^~(+{2{{4{(-2'sd0)}}}}));
  localparam signed [3:0] p15 = ((((-2'sd0)<(5'sd14))!=((4'd3)<<<(-4'sd3)))<(((-4'sd6)+(-2'sd1))&((2'd2)<<(2'd1))));
  localparam signed [4:0] p16 = ((((4'sd7)%(4'd13))<((-2'sd0)?(2'd0):(-5'sd15)))<=(((5'd13)?(2'd0):(2'd3))?((5'd9)?(3'sd1):(2'd2)):((-3'sd3)===(5'sd8))));
  localparam signed [5:0] p17 = {3{((-(5'd21))^(!(4'd8)))}};

  assign y0 = (((p4?a2:p2)!={4{p7}}));
  assign y1 = (|({(p7?b1:a2),(b3?a5:a4)}?((+a2)|(b0)):((a3)^~(b5))));
  assign y2 = (b3|b1);
  assign y3 = (~|(|((!(^b0))*(!(a2+a0)))));
  assign y4 = ({a1}?{p3,a5}:(a1&p4));
  assign y5 = (|($signed((|$unsigned($unsigned((~|{4{{2{a3}}}})))))));
  assign y6 = (!{(^b4),(p8<<p16)});
  assign y7 = ((a4?a3:b1)?(!(a3?a4:p13)):(p14?a4:a0));
  assign y8 = (4'd13);
  assign y9 = ((^(b2?p3:a1))?(&$signed(p4)):(~&(~|p3)));
  assign y10 = (((p0<a3)?(b4?p10:a4):(~^(-5'sd15)))^($unsigned((5'sd3))^((2'd2)^(b1<<p15))));
  assign y11 = (|((~(p17||p3))/p2));
  assign y12 = (+((2'd1)<<<{2{p7}}));
  assign y13 = (2'sd0);
  assign y14 = ((b0^p16)/b3);
  assign y15 = ((4'd2 * (b2||b0))^~(^(^($signed((a1^~a0))!==((b5*b0))))));
  assign y16 = ({2{({2{a3}}|{2{b2}})}}>(({2{a5}}===(b1^~a2))!=={2{{3{b3}}}}));
  assign y17 = {(-{p15}),(^(p9<p11)),(3'd6)};
endmodule
