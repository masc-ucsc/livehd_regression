module expression_00861(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd2 * ((3'd2)||(2'd0)));
  localparam [4:0] p1 = (~|(4'd11));
  localparam [5:0] p2 = ((|((4'd3)>=(-4'sd0)))<<<((3'd0)<=(-5'sd4)));
  localparam signed [3:0] p3 = (^(2'sd1));
  localparam signed [4:0] p4 = {((-3'sd3)&(3'd2)),{(3'sd1),(3'd5),(-2'sd1)}};
  localparam signed [5:0] p5 = (|((-(&(&((5'd21)===(-4'sd0)))))^({2{(4'd0)}}>=((4'd4)?(2'd2):(2'd2)))));
  localparam [3:0] p6 = {(((5'd17)?(2'sd0):(2'd0))?((4'd7)?(3'd3):(5'd0)):{(5'd9),(5'd17),(4'd10)}),(2'sd0)};
  localparam [4:0] p7 = ((5'd11)!==(4'd4));
  localparam [5:0] p8 = (6'd2 * (!(-(5'd12))));
  localparam signed [3:0] p9 = ((-2'sd0)*((5'd5)&&(-5'sd14)));
  localparam signed [4:0] p10 = (((3'd1)<<(3'd2))+(+(-4'sd7)));
  localparam signed [5:0] p11 = (+{{((-3'sd0)-(3'd1)),(!(|(2'd0)))},(!((-(!(5'd27)))<<<((4'sd5)==(2'sd1))))});
  localparam [3:0] p12 = ((3'd5)<<(4'sd3));
  localparam [4:0] p13 = (((|(3'd3))&&((3'd0)?(4'sd6):(2'd2)))!==(((4'sd5)-(5'sd13))?((-4'sd4)?(2'd3):(3'd5)):(~^(5'd23))));
  localparam [5:0] p14 = (((-5'sd10)%(-5'sd2))>>((4'd11)/(5'd4)));
  localparam signed [3:0] p15 = {3{((5'd15)<<(3'd5))}};
  localparam signed [4:0] p16 = ({4{(2'd0)}}!=((4'd15)-(3'sd1)));
  localparam signed [5:0] p17 = (~((((-2'sd1)>(2'd2))!={((3'd1)&(2'sd0))})===(2'sd1)));

  assign y0 = (p11?b5:p1);
  assign y1 = (a2?a4:b5);
  assign y2 = (~|$signed($unsigned((5'd2 * p0))));
  assign y3 = {{p5,b1,a0},(-b5),(&a0)};
  assign y4 = {1{{4{p10}}}};
  assign y5 = {(~^p6),(|b3)};
  assign y6 = ({3{{1{(p16)}}}});
  assign y7 = {(3'd2),(~(5'd23)),(4'd13)};
  assign y8 = $signed($signed($signed($unsigned((($unsigned((~&a2))?((+b2)):((^b3))))))));
  assign y9 = (~^{4{(p9-p9)}});
  assign y10 = {3{{{3{a3}},{p5,p13}}}};
  assign y11 = ((^(p13>>>p6))|(~^(5'd2 * b0)));
  assign y12 = ((a4?p6:p10)?{1{(!a5)}}:(~(p12>>>p7)));
  assign y13 = (|(|{(|a4),(-p2),{a4}}));
  assign y14 = (~^((^$unsigned(p16))%p0));
  assign y15 = (~(!{({(b2-p1),(p0?p11:p0)}>(4'd5))}));
  assign y16 = ({b2,p8,b5}?{a1,p0}:(+(p17<=p12)));
  assign y17 = $signed((2'd0));
endmodule
