module expression_00558(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({3{{1{(4'd12)}}}}?({1{(-5'sd12)}}>=(-(5'sd5))):({(3'sd2)}>((5'sd12)||(-3'sd1))));
  localparam [4:0] p1 = {(!((4'd13)?(-5'sd6):(3'sd0))),((4'd13)?(3'd0):(-4'sd4)),((5'd2)?(2'sd0):(3'd3))};
  localparam [5:0] p2 = (((4'sd6)^(-4'sd4))?(|(4'sd4)):{3{(2'sd0)}});
  localparam signed [3:0] p3 = (&(4'sd3));
  localparam signed [4:0] p4 = ((((5'd30)||(5'd2))>>((4'd10)-(4'd13)))<=(((5'd17)^~(5'sd7))&&((5'd16)>(3'sd1))));
  localparam signed [5:0] p5 = (((-3'sd1)^~(2'd3))|(-2'sd1));
  localparam [3:0] p6 = ((4'd11)?(3'd6):(-2'sd0));
  localparam [4:0] p7 = ((5'd20)===((-4'sd6)?(-2'sd1):(3'sd1)));
  localparam [5:0] p8 = ((+(((-4'sd6)?(-3'sd2):(-3'sd0))===(-(~^(5'sd11)))))>=((~(5'd26))?((-3'sd2)?(-4'sd1):(5'd17)):((5'sd4)?(5'sd8):(4'sd7))));
  localparam signed [3:0] p9 = ((5'd22)?(4'sd6):(~|((5'sd0)==(2'sd0))));
  localparam signed [4:0] p10 = {4{((-2'sd0)+(3'd2))}};
  localparam signed [5:0] p11 = (^(^((~|{(-3'sd3)})<=(-{(2'd2)}))));
  localparam [3:0] p12 = (~^(6'd2 * (3'd1)));
  localparam [4:0] p13 = (((5'sd8)|(2'sd1))%(3'sd0));
  localparam [5:0] p14 = {2{({(5'd27),(2'sd1)}<<<(4'd2 * (4'd12)))}};
  localparam signed [3:0] p15 = ({((-3'sd0)|(3'sd0)),((3'sd0)>(4'sd7)),(+((2'd2)&&(2'sd1)))}&&{(~|((2'd1)<<(2'd1))),{2{(+(3'd7))}}});
  localparam signed [4:0] p16 = (~|(3'd0));
  localparam signed [5:0] p17 = {3{(~^(2'd2))}};

  assign y0 = ((4'd2 * (p0&a1))!={4{b1}});
  assign y1 = (~((3'd0)?(~(5'd22)):(-5'sd8)));
  assign y2 = (~&(~((+((a0!=p17)>=(-b2)))&&((^p10)?(a0-a3):{3{b5}}))));
  assign y3 = (2'sd1);
  assign y4 = (((~|$signed(p9))*(^(~|b0))));
  assign y5 = (~^(!(|{(|(|{3{p10}})),{a2,p8,a4},(&{4{p9}})})));
  assign y6 = (4'sd1);
  assign y7 = (&((~b1)?(p12?p8:p8):(a0?p10:p15)));
  assign y8 = ($signed($signed(a0))===$signed((a0>b0)));
  assign y9 = (b1<<a3);
  assign y10 = $signed(((({1{b2}}<$unsigned(p11))^{2{{4{a4}}}})>>$unsigned($signed((($signed({3{a2}})<<(b3|a0)))))));
  assign y11 = $unsigned({{b0},(b2>=a0)});
  assign y12 = (+$signed((~&(|($unsigned((&$signed($unsigned((!(+b3)))))))))));
  assign y13 = (+{4{(p11<<<p16)}});
  assign y14 = (~{(+{((~&(p12<<p12))<<<(4'd10))}),((4'd7)<(-(|(p15>>p2))))});
  assign y15 = (4'sd2);
  assign y16 = (a2>>p14);
  assign y17 = (+$unsigned(p9));
endmodule
