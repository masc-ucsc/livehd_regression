module expression_00794(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd26);
  localparam [4:0] p1 = (~&({1{({1{(5'd21)}}?((-2'sd0)>=(3'sd2)):((4'd8)?(3'sd0):(4'd14)))}}+(^(|(((5'd24)?(-4'sd2):(4'd8))=={1{(2'sd0)}})))));
  localparam [5:0] p2 = {((5'sd3)?(3'sd2):(5'sd10)),((~|(3'd3))-((4'sd5)|(4'sd2))),{(3'sd1),(-4'sd2),(-2'sd0)}};
  localparam signed [3:0] p3 = ((&(^((-4'sd6)===(4'd12))))<=((3'd3)?(3'd2):(2'd3)));
  localparam signed [4:0] p4 = ((|{((5'd18)<<(-5'sd7)),{(-2'sd1),(4'sd7),(5'd1)}})==(!(-({(5'd21),(5'd16),(-3'sd1)}+{(4'sd3),(3'd2),(3'd1)}))));
  localparam signed [5:0] p5 = ({(5'd5),(5'd14)}?(&(4'd3)):((4'sd7)?(-5'sd9):(-3'sd2)));
  localparam [3:0] p6 = (5'd13);
  localparam [4:0] p7 = (!{4{(((-4'sd0)||(2'sd1))>>>{3{(5'd21)}})}});
  localparam [5:0] p8 = {(+(+(((2'sd0)-(5'd8))&&(~^(3'd1))))),(~&((-(6'd2 * (4'd3)))&&((2'd1)&(-2'sd1))))};
  localparam signed [3:0] p9 = ({4{((3'sd1)===(3'd5))}}+(((3'd7)!==(5'sd9))|{3{(4'd1)}}));
  localparam signed [4:0] p10 = (((2'd1)+(5'sd11))+((3'sd3)>>(3'sd2)));
  localparam signed [5:0] p11 = (^(((!(-4'sd6))|((5'd6)?(-3'sd3):(-4'sd7)))>((6'd2 * (4'd12))?((3'd4)!=(5'd2)):((5'sd4)?(4'd5):(-5'sd11)))));
  localparam [3:0] p12 = ({{3{(2'd2)}}}<<{((5'd6)|(-3'sd2)),((5'sd15)<<(4'd5)),((2'sd0)|(-4'sd0))});
  localparam [4:0] p13 = (&(2'd2));
  localparam [5:0] p14 = ({4{(5'sd11)}}?{(4'sd4),(2'd2),(5'd3)}:{(-4'sd1),(-3'sd0)});
  localparam signed [3:0] p15 = (!((!(-((-3'sd0)?(2'd1):(-4'sd0))))>(&((4'sd7)?(4'd4):(3'sd0)))));
  localparam signed [4:0] p16 = {{1{(3'd2)}},((5'sd14)&&(2'sd1)),((4'sd6)==(2'd0))};
  localparam signed [5:0] p17 = (~&(|(+(&{(~&(~{2{{(-2'sd0),(5'd2)}}}))}))));

  assign y0 = (-5'sd12);
  assign y1 = ((2'd3)>(5'd1));
  assign y2 = (a0?a1:p4);
  assign y3 = (((p4?p6:p16)?(p4?a4:p1):(p4?p8:a1))|((6'd2 * p0)?(a5!==a2):(p5)));
  assign y4 = (b2===b4);
  assign y5 = (+((!(~|p2))?(-(p3?p2:p5)):(5'd27)));
  assign y6 = (~^(~&(-2'sd0)));
  assign y7 = (-3'sd1);
  assign y8 = $unsigned($unsigned((3'd0)));
  assign y9 = $signed({3{{p17,p12,p5}}});
  assign y10 = (((|({1{(b4)}}))?((b4<=a1)>$signed(a3)):((^p3)+$signed(a5))));
  assign y11 = {2{(|({2{b0}}&{3{a2}}))}};
  assign y12 = ((&(p7^p16)));
  assign y13 = $signed((2'd3));
  assign y14 = {2{a4}};
  assign y15 = ((-a5)<<<(a1?a5:b2));
  assign y16 = (((&(-$signed(p8)))==((p8<=p10)))&&$unsigned(($signed({2{p2}})>(p12||p7))));
  assign y17 = (4'd7);
endmodule
