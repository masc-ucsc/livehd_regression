module expression_00432(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(2'd1));
  localparam [4:0] p1 = (4'd11);
  localparam [5:0] p2 = ((((3'd1)?(-3'sd3):(3'd4))==((-5'sd10)&&(5'd21)))<<<(((2'd3)?(-5'sd1):(3'd0))!=((4'd14)>(2'd3))));
  localparam signed [3:0] p3 = (+(4'sd2));
  localparam signed [4:0] p4 = ((~(((-2'sd1)&(4'd8))<((-5'sd7)>=(5'd20))))||(((4'd4)%(2'sd0))+(~|((5'd13)?(3'sd0):(3'sd1)))));
  localparam signed [5:0] p5 = {{2{({(5'sd9),(2'sd0)}<<((5'd9)-(-2'sd1)))}},{3{{4{(5'sd3)}}}}};
  localparam [3:0] p6 = (-5'sd5);
  localparam [4:0] p7 = ({1{(3'd6)}}?(5'd16):{1{((5'd10)?(5'd0):(3'd1))}});
  localparam [5:0] p8 = (4'd10);
  localparam signed [3:0] p9 = {{(-3'sd1),(-5'sd13)},((2'sd1)^(5'd12)),((4'sd0)?(2'd3):(5'sd7))};
  localparam signed [4:0] p10 = ({4{(2'sd1)}}!=={1{(2'sd1)}});
  localparam signed [5:0] p11 = {(((3'sd2)?(2'd2):(-3'sd2))|(&(+(2'd3)))),(+(((3'sd2)?(-4'sd2):(-5'sd7))>>>(-(4'sd1))))};
  localparam [3:0] p12 = ((((2'd2)+(4'd5))!==(5'd2 * (5'd21)))?(((-5'sd15)|(4'd2))<<(^(2'd1))):{(2'sd0),(4'sd7),(3'sd0)});
  localparam [4:0] p13 = ((((3'd6)<<(2'sd1))<((4'd5)===(4'd0)))<<<(^(-{2{(-2'sd0)}})));
  localparam [5:0] p14 = (+(((~&(+(-3'sd3)))^(!(+(4'd6))))!=(5'd2 * (&(|(2'd0))))));
  localparam signed [3:0] p15 = (~(((+(-3'sd1))<((-4'sd2)||(2'sd1)))-(((3'd7)<(5'd14))^~{2{(2'd0)}})));
  localparam signed [4:0] p16 = (5'd12);
  localparam signed [5:0] p17 = (-{(^((-3'sd2)|(4'd15))),{{(2'sd1)},((-3'sd0)>=(4'd13))}});

  assign y0 = $unsigned((4'sd2));
  assign y1 = {2{(-5'sd12)}};
  assign y2 = ((|(p8%p3))>=(a0^p5));
  assign y3 = ((~{2{b2}})?(b4?a1:a0):{4{b0}});
  assign y4 = (5'd22);
  assign y5 = (4'd15);
  assign y6 = (p16&a2);
  assign y7 = {2{(|(4'sd1))}};
  assign y8 = ((~^{3{{b1,p17}}})+{(-4'sd5)});
  assign y9 = (~|{2{a5}});
  assign y10 = (^(-(~(|(!(~^(!(^(~|{1{(!{2{a4}})}})))))))));
  assign y11 = (~&{1{{2{((b2?b2:b3)?(p11?a4:a1):(~&b2))}}}});
  assign y12 = {1{((!(~&(~|(b0<<a3))))===((b4|b4)!=(a3^b2)))}};
  assign y13 = ((&(p12?b3:p16))?(|(p9?b2:b3)):(p10?p10:a5));
  assign y14 = {4{{3{(~b5)}}}};
  assign y15 = {4{{3{a3}}}};
  assign y16 = ({3{(p11>>>p15)}}||(((p13>>p11)||{3{p0}})&{1{(p12^~p9)}}));
  assign y17 = (~|($signed($unsigned(($unsigned(a4)?(b5===a5):(~p11))))&($signed(((p1^~b5)<=(a2?b0:b4))))));
endmodule
