module expression_00210(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(&{4{(3'd4)}}));
  localparam [4:0] p1 = (|(-5'sd11));
  localparam [5:0] p2 = ((2'd3)?(4'd1):(5'sd5));
  localparam signed [3:0] p3 = ((2'd3)?(((4'd1)!=(-4'sd2))&((2'd0)>>>(5'sd11))):{4{(2'd1)}});
  localparam signed [4:0] p4 = (((2'd3)&(-3'sd3))==(-(6'd2 * (2'd1))));
  localparam signed [5:0] p5 = (2'd2);
  localparam [3:0] p6 = (~&(((-2'sd0)?(2'd0):(-4'sd5))?(!(5'sd4)):(&(2'd1))));
  localparam [4:0] p7 = (4'sd5);
  localparam [5:0] p8 = (|(5'd27));
  localparam signed [3:0] p9 = {1{(|(2'd2))}};
  localparam signed [4:0] p10 = (|(((3'd2)*(4'd11))&&((4'd6)==(-3'sd1))));
  localparam signed [5:0] p11 = (5'd2);
  localparam [3:0] p12 = ((((2'd1)?(2'd2):(-4'sd6))?(3'd2):((2'sd1)&(3'd1)))^~(((|(-5'sd13))-((4'd10)+(-2'sd1)))!=((3'd6)?(5'd8):(-2'sd1))));
  localparam [4:0] p13 = {{(-((-3'sd3)^(3'sd1))),{(4'sd1),(3'sd0)},(+((-5'sd7)?(5'd26):(3'd0)))},((2'd1)|(~(+((4'd6)===(2'd0)))))};
  localparam [5:0] p14 = ((~|(5'd10))==(5'd7));
  localparam signed [3:0] p15 = ((((2'd1)<<(4'sd1))!==((3'd5)!=(4'sd7)))>>>(!((-4'sd1)>>>(4'sd1))));
  localparam signed [4:0] p16 = (4'd5);
  localparam signed [5:0] p17 = (2'd0);

  assign y0 = ((p6>p13)?(p16?p13:p1):(p10?p9:p0));
  assign y1 = (~&{(&p11),(!b5)});
  assign y2 = ({4{p17}}<<<(^{2{p16}}));
  assign y3 = (~({3{(b0>>>b3)}}^~(-{4{(a4!==b5)}})));
  assign y4 = {({(a1<<b1),(!b0)}-((|a5)|(~&p0))),(((a2)>=(a4&a4))>=((^b5)!==(~&b4)))};
  assign y5 = (((a3!==a5)&&(b4!=p12))>((b2>>p2)?(b0<<a3):(a5>>>a3)));
  assign y6 = (2'd0);
  assign y7 = (((a4===b5)==(a0|b0))>((b5!==a0)!=(-2'sd1)));
  assign y8 = (((p10+b5)^(p13?b0:p6))?((4'd2 * b1)?(p15<<p13):$unsigned(p3)):$unsigned(((b4||p8)+(b1>b1))));
  assign y9 = (^(2'd2));
  assign y10 = (($signed((&b5))!={3{b2}})<(~({4{a0}}!==(b4<b1))));
  assign y11 = ((a2?b2:b4)%b1);
  assign y12 = $unsigned($signed(({(p16?p16:p14),(p15),(p5?p9:p2)}?$signed((~&{(~^p15)})):(3'd4))));
  assign y13 = {4{{2{b2}}}};
  assign y14 = (6'd2 * {b0,b2});
  assign y15 = (-4'sd0);
  assign y16 = ((+(&(!(b4===b0))))<(3'd4));
  assign y17 = $signed(((a5<<b5)===(b0!==a4)));
endmodule
