module expression_00814(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~({4{(-4'sd3)}}!==((2'sd1)>(3'sd0))));
  localparam [4:0] p1 = ((((2'sd0)<<<(-2'sd1))||(|(5'sd0)))===(^((-4'sd5)&&(5'sd15))));
  localparam [5:0] p2 = ((~(-5'sd2))>>(5'sd7));
  localparam signed [3:0] p3 = (3'sd3);
  localparam signed [4:0] p4 = (({(5'd2 * (4'd12))}!==((6'd2 * (2'd1))-{(4'd0)}))-({{((2'sd1)===(-4'sd6))}}+(!(!(!(-4'sd1))))));
  localparam signed [5:0] p5 = (({(-4'sd4),(-3'sd2)}<<{1{(-4'sd2)}})!==(5'd10));
  localparam [3:0] p6 = (~(((-(3'd6))<((2'sd1)?(3'd4):(2'sd1)))?(~|((2'sd1)?(2'd3):(4'd10))):(~^(~|((4'd10)&(2'd3))))));
  localparam [4:0] p7 = ({(-3'sd0),(-3'sd2),(-5'sd13)}?((-4'sd4)?(2'sd1):(3'd0)):{(5'd20),(4'd7)});
  localparam [5:0] p8 = {2{{4{(5'sd6)}}}};
  localparam signed [3:0] p9 = (&({((5'sd0)<<<(3'd3)),((-3'sd0)^(5'd30))}?(&{2{((5'd20)?(-4'sd6):(2'd1))}}):((+(2'd0))?(^(2'sd0)):(+(3'd4)))));
  localparam signed [4:0] p10 = (-2'sd1);
  localparam signed [5:0] p11 = ((((-2'sd0)^~(3'd3))?((-4'sd1)?(3'd1):(3'd0)):((2'd2)?(2'd2):(4'd4)))!==(((-3'sd0)<(-4'sd0))!==(~((5'd18)?(4'd15):(-3'sd2)))));
  localparam [3:0] p12 = (~|(3'd7));
  localparam [4:0] p13 = (~&(~&((((5'd30)==(3'd6))===(!(4'd5)))>>(~((5'sd13)!==(5'sd2))))));
  localparam [5:0] p14 = (^(((~^(3'd6))?((3'sd3)-(2'sd0)):((4'sd7)?(3'd1):(5'sd11)))?((+(2'd1))?((2'sd1)?(4'sd4):(-2'sd1)):((-3'sd0)==(4'd9))):((5'd29)?(&(-2'sd1)):(3'sd1))));
  localparam signed [3:0] p15 = (((((-5'sd14)<<<(3'sd2))>>((2'd2)===(-5'sd7)))!==((4'd2 * (3'd0))===((2'd1)<<<(4'sd3))))!==((((-4'sd2)<=(2'd1))<<((5'sd1)!=(4'd3)))<=(((5'd1)>>(3'd3))&&((5'd31)<(-5'sd13)))));
  localparam signed [4:0] p16 = (~&((!((~^(5'd0))?(~(-3'sd3)):((2'sd0)!==(5'd17))))<<<{3{{1{(4'd9)}}}}));
  localparam signed [5:0] p17 = {({(3'd0),(3'sd2),(5'sd4)}?{((4'sd5)>>(4'd1))}:((3'sd0)?(5'd21):(5'd27)))};

  assign y0 = ($signed((-((~&b3)<(~^b5))))<<{({a1,a5,b5}&&{4{a3}})});
  assign y1 = (((a3!=a4)|{1{{3{b0}}}})+({1{{3{a1}}}}!==(a2<=a1)));
  assign y2 = {{(p4?p2:p1),((5'd8)+{p14,p15})},{3{(3'd1)}}};
  assign y3 = (((p1-b4)<=(a2%p2))-((|(p10))^~(^(4'd2 * p12))));
  assign y4 = (((~(b3?a2:a5))!=$signed((a0?b3:a2)))&&(|((+$unsigned((b2?b1:a3)))^{4{b1}})));
  assign y5 = {{(a5|b2)},{p10,p11,p13}};
  assign y6 = (-(4'd2 * (a2<p1)));
  assign y7 = {1{({(b1?p12:p10),$signed(p5)}?{(p17?b1:p16)}:{1{(p4?p5:a1)}})}};
  assign y8 = {4{$unsigned((p0<p8))}};
  assign y9 = (3'd3);
  assign y10 = (((p16&&b1)?(p11?p9:p11):(p8<p9))<<((-p1)?(-p13):(-p17)));
  assign y11 = (-(~&((-4'sd1)-(~(4'sd2)))));
  assign y12 = (($unsigned((2'd3))<<<(4'd7))^~(((4'd5)?(b1>b5):(2'd2))==(3'sd3)));
  assign y13 = ((5'd2 * a0)-(a3));
  assign y14 = (~|((!(b1?b3:a3))!==((a4==a5)!==(a0<<<b1))));
  assign y15 = (((p15?a0:p5)>>>((p17<<p1)&&(b3||a3)))<<((-3'sd3)<(2'sd0)));
  assign y16 = {1{{3{(b4?p3:p13)}}}};
  assign y17 = $unsigned(($signed(((p1?p8:p8)?(p5?p6:p4):(p8?p1:p2)))?$signed(((p1?p12:a5)?$signed(p11):(p8?p9:p14))):(((a1?b4:p7)?(p1?b5:p17):(p5|p8)))));
endmodule
