module expression_00341(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(^(~|{1{{3{(-4'sd5)}}}})));
  localparam [4:0] p1 = {(((4'd15)>(3'd0))!==((4'sd1)!=(5'd9))),({(2'd0),(-4'sd1)}|(~{(-5'sd4)}))};
  localparam [5:0] p2 = ((6'd2 * ((4'd7)^~(4'd7)))===(((4'd6)||(-2'sd1))<=(~^{2{(-4'sd0)}})));
  localparam signed [3:0] p3 = (({4{(4'sd4)}}===((-5'sd5)<<<(2'sd0)))^~({4{(-2'sd0)}}?((2'd3)?(2'sd1):(5'sd3)):{1{(3'sd2)}}));
  localparam signed [4:0] p4 = ({2{((3'sd3)^(3'sd3))}}>{1{((-5'sd6)|(-3'sd3))}});
  localparam signed [5:0] p5 = ({(4'd0)}!={(5'sd2),(4'd14)});
  localparam [3:0] p6 = ((~&{(|(5'd29))})-((5'sd5)?(4'd12):(-3'sd2)));
  localparam [4:0] p7 = (^(((3'd3)&(-2'sd1))*(~&(+(-2'sd1)))));
  localparam [5:0] p8 = (~|(^((2'd3)<(4'd4))));
  localparam signed [3:0] p9 = (4'd15);
  localparam signed [4:0] p10 = ((((-2'sd0)>(-4'sd0))?((4'sd7)?(-5'sd13):(3'd5)):((3'sd0)==(4'd2)))!=(((-5'sd14)?(3'd7):(2'd0))?((4'd15)?(3'd6):(4'sd6)):((5'd30)+(3'sd0))));
  localparam signed [5:0] p11 = ((5'd29)?(4'd13):(3'd7));
  localparam [3:0] p12 = {2{{1{(-4'sd0)}}}};
  localparam [4:0] p13 = (6'd2 * ((3'd0)?(2'd1):(2'd2)));
  localparam [5:0] p14 = {{{4{(4'd6)}},{(2'sd0),(4'd2)}},(~{4{(-3'sd3)}})};
  localparam signed [3:0] p15 = (((4'd15)%(5'sd12))%(3'sd3));
  localparam signed [4:0] p16 = ((4'sd2)?(-4'sd3):(-4'sd7));
  localparam signed [5:0] p17 = {3{{4{(5'd16)}}}};

  assign y0 = {{p17,p8,b4}};
  assign y1 = $unsigned(p15);
  assign y2 = (!(~(-3'sd2)));
  assign y3 = (((~$unsigned(a3))&$unsigned((a1|p6))));
  assign y4 = $signed((((p16&&p2)%b5)+((p5|a0)>$unsigned((p15<=b3)))));
  assign y5 = (!$unsigned($unsigned(((p13<<<b0)|{b1,p2}))));
  assign y6 = (~&(2'd1));
  assign y7 = ((~^(b0!==b5))<<({b3,b5}>$signed(b0)));
  assign y8 = {1{({2{{2{{1{p13}}}}}}>(&{4{{2{b0}}}}))}};
  assign y9 = (^((|(b4?p13:b0))?(3'd4):{1{((-3'sd2)>=(b4?p13:p0))}}));
  assign y10 = (4'd2 * (b0?b0:p0));
  assign y11 = (~&{{(&((!b4)?(&a5):(+a3)))},{{(b1?b3:b1)},{a0,a2,a3},{(-a3)}}});
  assign y12 = (!{{1{$unsigned((|{1{p5}}))}}});
  assign y13 = {{b4}};
  assign y14 = {1{(({1{{2{(b5>>a2)}}}}?(-3'sd0):((+(b3?a2:a4))==(a5<<a5))))}};
  assign y15 = ((p12^~p6)|(a0>>a2));
  assign y16 = $unsigned({1{(!{({p6}^(!b2)),{{1{b4}},{3{b0}},{b5,p9}},((|a5)^{2{a1}})})}});
  assign y17 = (+(^{1{(|p4)}}));
endmodule
