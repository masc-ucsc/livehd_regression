module expression_00131(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-{2{(-2'sd1)}})?(2'd2):((2'd2)?(4'sd3):(3'sd2)));
  localparam [4:0] p1 = (-(-4'sd2));
  localparam [5:0] p2 = (-3'sd1);
  localparam signed [3:0] p3 = (-({1{(2'd2)}}?((-2'sd1)?(3'sd2):(-2'sd0)):((4'sd1)&&(3'd2))));
  localparam signed [4:0] p4 = {({((-4'sd2)^(4'd8))}||((-5'sd3)!=(2'd2)))};
  localparam signed [5:0] p5 = (&((((2'd3)||(5'd11))&&{(5'd28),(5'd12)})&&(((-2'sd0)!=(5'd22))>((3'd7)+(-5'sd14)))));
  localparam [3:0] p6 = ((((4'd3)&&(4'd1))?((2'd2)^(2'd3)):((5'd2)?(4'sd0):(3'sd1)))>>(((2'd0)>=(-2'sd1))?((-5'sd15)/(4'd8)):((-2'sd0)?(5'sd0):(3'd1))));
  localparam [4:0] p7 = ((-5'sd9)<<(4'sd5));
  localparam [5:0] p8 = {4{((3'd7)===(3'd2))}};
  localparam signed [3:0] p9 = ((((3'd5)!=(-2'sd0))<(6'd2 * (2'd3)))?((~(4'd2))==((5'sd10)===(2'd1))):({(5'd19),(5'd6)}!=((-5'sd14)>>>(5'sd9))));
  localparam signed [4:0] p10 = ((((-5'sd2)?(5'd24):(4'sd2))?((-3'sd3)?(5'sd3):(5'sd2)):(2'sd1))^(((3'sd2)||(2'd3))?((5'd22)|(-5'sd6)):(2'sd0)));
  localparam signed [5:0] p11 = ((!((4'd13)?(2'd1):(2'd1)))?(&(!((2'd0)?(5'sd2):(-3'sd3)))):((-(3'sd3))?(|(-2'sd1)):(-(4'd13))));
  localparam [3:0] p12 = ((+(-4'sd0))<(((5'd13)>=(5'd25))|{4{(3'd3)}}));
  localparam [4:0] p13 = {4{(~(2'sd1))}};
  localparam [5:0] p14 = (+(~(((5'sd1)?(-4'sd3):(-3'sd0))<<<((5'd15)!=(5'sd1)))));
  localparam signed [3:0] p15 = ({(3'd3),(2'sd1),(5'sd14)}?({(2'd3)}>>((-2'sd1)&&(-5'sd7))):{(~&(5'd21)),(~^(2'd2))});
  localparam signed [4:0] p16 = {1{(~&((~&(+(+(5'd22))))<={(2'sd0),(-3'sd2),(4'd13)}))}};
  localparam signed [5:0] p17 = ((((3'sd0)?(2'd3):(3'd2))?((5'd22)?(5'd16):(-5'sd1)):((-5'sd7)?(3'sd3):(5'sd1)))?(((-2'sd0)?(3'd6):(3'd0))?((3'sd2)?(2'sd0):(-3'sd1)):((2'd0)?(4'sd5):(3'sd2))):(((2'd2)?(3'sd1):(2'd2))?((-4'sd4)?(-5'sd2):(4'd9)):((-2'sd1)?(3'sd2):(5'd0))));

  assign y0 = {{3{{{4{p7}},{p12,p10},{4{p7}}}}}};
  assign y1 = (-5'sd13);
  assign y2 = {{2{p4}},((a5?b3:a5)),(a4?b3:p3)};
  assign y3 = {({2{p6}}-{2{p7}}),(~{1{{3{p8}}}}),{(p13+p11),(+p15),(p8!=p8)}};
  assign y4 = (((p17?p13:p4)>=(a3?p15:p11))?(~(^((+a5)<<(^p1)))):(&(!((p8?p16:p17)?(~^p7):(p1?p12:p11)))));
  assign y5 = (&({4{a2}}+((a4==b0)===$signed(a2))));
  assign y6 = (|(~|(~|(~^(~^a0)))));
  assign y7 = {1{{2{{3{a0}}}}}};
  assign y8 = (+{3{p6}});
  assign y9 = (~|(~|(~|(-(|(!(-(&(~|(~(~^(~(^(~|(!(~&p16))))))))))))))));
  assign y10 = ((&((a4===a2)?(b2?a0:a5):(&a5)))?(^((b3!=b4)>=(b2?b0:b5))):(!((~^a1)>>>(b4/b1))));
  assign y11 = ((~|((|b2)==(|b2)))&(+((a4&a5)>$unsigned(a4))));
  assign y12 = (4'd12);
  assign y13 = ({1{{1{(({4{a4}}|(a4>>>b2))||({4{b5}}===((b3>>b5))))}}}});
  assign y14 = ((p13?p7:p6)>((p4?p5:p1)|(p13?p11:p4)));
  assign y15 = (((b3?p4:a3)?(a3?b3:p15):(|{3{a0}}))<{2{(p16?b1:b0)}});
  assign y16 = (-((5'd14)?(&{a0,a3,a0}):{(+a5)}));
  assign y17 = {4{((p8?p1:p5)|(2'd2))}};
endmodule
