module expression_00752(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd1),(4'd1),(-5'sd15)};
  localparam [4:0] p1 = (|(((&(-3'sd1))<<((-4'sd4)==(5'd21)))&((+(-2'sd0))&&((3'd6)^(-4'sd6)))));
  localparam [5:0] p2 = ((3'sd0)?(4'sd3):(-3'sd2));
  localparam signed [3:0] p3 = (-4'sd0);
  localparam signed [4:0] p4 = ((4'sd0)?{2{(4'sd3)}}:{2{(-3'sd2)}});
  localparam signed [5:0] p5 = (2'sd1);
  localparam [3:0] p6 = (((5'd30)?(5'd8):(-5'sd15))?{(2'd3),(5'sd1),(4'd8)}:{4{(4'd0)}});
  localparam [4:0] p7 = (5'd2 * (5'd11));
  localparam [5:0] p8 = (({1{(-5'sd6)}}!=((-5'sd1)-(-4'sd4)))!==(((2'sd0)===(-5'sd0))^((5'sd13)&(4'd5))));
  localparam signed [3:0] p9 = (~(&(3'd0)));
  localparam signed [4:0] p10 = (&((((4'd9)?(4'd3):(4'sd4))+{3{(-3'sd0)}})<<<((4'sd7)?(3'd5):(4'd9))));
  localparam signed [5:0] p11 = (((5'd9)<<((2'd2)<=(-4'sd6)))?((2'sd0)?(-3'sd1):(2'sd0)):(~&((2'd3)-(3'sd3))));
  localparam [3:0] p12 = (4'd15);
  localparam [4:0] p13 = ({3{{(3'd4),(-3'sd2),(-3'sd2)}}}=={((5'd26)?(-5'sd15):(5'd6)),{(-4'sd4),(2'd0)}});
  localparam [5:0] p14 = (((-3'sd2)|(4'd1))?((4'd11)<<<(5'd9)):(-4'sd6));
  localparam signed [3:0] p15 = {2{(-5'sd9)}};
  localparam signed [4:0] p16 = ({4{(-3'sd2)}}?{(3'sd3),(-2'sd1),(-2'sd1)}:((-2'sd1)!=(2'sd1)));
  localparam signed [5:0] p17 = (((-2'sd0)?(3'sd1):(4'd7))%(2'sd1));

  assign y0 = $unsigned(p17);
  assign y1 = {4{(p15>>>p1)}};
  assign y2 = (~&((~&(~&(a5+p6)))<<<(|$unsigned((p6^p12)))));
  assign y3 = (~(!(p11>>p12)));
  assign y4 = ($signed(a0)?(+p7):(4'd12));
  assign y5 = (|((p16|a1)>{2{p2}}));
  assign y6 = (({3{b3}}&&{4{b4}})==({3{p7}}<{1{(a4<<<p2)}}));
  assign y7 = {p10,p17};
  assign y8 = {(p13&p0),(p13?p13:p16),{2{b5}}};
  assign y9 = (2'sd0);
  assign y10 = (((6'd2 * (p6||p1))-{(5'd2 * p6),{p12,p4}})+({(a0!==a2)}+((~^b4)&(-p13))));
  assign y11 = {({((p5^~p1)?(|(p4>>p1)):{p1,p1,p2})}>>>({(p0?p0:p0)}&{(p10|p7),(p4||p8),(p14<<<p9)}))};
  assign y12 = (((b3+p11)<<{a3,b1})?{(&(b0&p8)),(a4?b3:a1)}:((b3?a1:b3)|{b0,b1}));
  assign y13 = (~^{2{(5'sd11)}});
  assign y14 = (~^{({p5,p11}>>>(^p9)),(+{a1,p15,p11})});
  assign y15 = (~((b5?a2:a5)?(b5?a3:b2):(a5?a1:b5)));
  assign y16 = (^$unsigned((((p16))^~(a5?p9:a4))));
  assign y17 = {4{(~&(a4<<<a4))}};
endmodule
