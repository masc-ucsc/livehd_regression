module expression_00890(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(|({3{(3'd5)}}!=((-3'sd2)!=(3'd4))))}};
  localparam [4:0] p1 = {1{(|(((2'sd0)?(-2'sd1):(5'd27))?((3'sd0)?(5'd22):(3'd4)):((-3'sd1)&(5'd12))))}};
  localparam [5:0] p2 = (5'd2 * {(2'd1),(3'd3)});
  localparam signed [3:0] p3 = (-(2'sd1));
  localparam signed [4:0] p4 = ({3{{1{(3'd1)}}}}!={2{((2'd0)>=(-4'sd4))}});
  localparam signed [5:0] p5 = (|((-2'sd1)?(5'd31):(4'd3)));
  localparam [3:0] p6 = {3{(2'sd0)}};
  localparam [4:0] p7 = (&(-3'sd0));
  localparam [5:0] p8 = (-{3{{4{(4'd12)}}}});
  localparam signed [3:0] p9 = (~^(2'sd0));
  localparam signed [4:0] p10 = (!(|(!({(3'sd2),(4'sd2)}&((3'd4)?(-3'sd1):(-2'sd0))))));
  localparam signed [5:0] p11 = ((3'sd2)!=={(~((5'sd13)+(5'sd12))),(-4'sd2)});
  localparam [3:0] p12 = (-3'sd0);
  localparam [4:0] p13 = ({3{(-4'sd4)}}?((3'd5)?(4'sd7):(3'd2)):((4'd6)?(4'd4):(5'd28)));
  localparam [5:0] p14 = ((((~|(-3'sd1))^((4'd1)==(-5'sd14)))!=((-(-5'sd0))>(-(3'd2))))<=(&(((5'sd9)^(4'd3))<<(~&(~^(5'd26))))));
  localparam signed [3:0] p15 = (((5'sd7)>>(4'd3))==((-5'sd12)!=(2'd0)));
  localparam signed [4:0] p16 = (+(-{3{(~|(^(3'sd0)))}}));
  localparam signed [5:0] p17 = (((5'd24)||(-4'sd5))<<((5'd9)%(-2'sd0)));

  assign y0 = ((-3'sd0)>>>(a4>>>b4));
  assign y1 = ({(a3|a5),(b0>=b0),(p3<=p7)}>={{(4'd2 * p8)},{3{p5}},{a0,p16,a1}});
  assign y2 = ({{a2,a0,a1}}^{{4{b2}},(b4<<a3),(p4|b3)});
  assign y3 = (^(2'd0));
  assign y4 = (($unsigned(b4)?{a2}:(b1?b0:a0))&$signed({((!a5)!==$signed(b0))}));
  assign y5 = (((p5<<<p2)?(b3!==b1):$signed(p7))?((a1===a2)?(p7?p11:p9):$unsigned(p2)):(((p14&&p1)&&$signed(p10))));
  assign y6 = {1{{2{{4{p2}}}}}};
  assign y7 = (5'd9);
  assign y8 = ((~(-2'sd1))-(~|{3{(b5^p7)}}));
  assign y9 = ((b3?b5:b0)^~(~^a2));
  assign y10 = (((6'd2 * b1)?{p15,p3,p15}:$signed(p8))?{(&{({b4,p9}&&(p5>=a0))})}:({p13,p15,p1}<$signed((b4?p14:p9))));
  assign y11 = (-4'sd1);
  assign y12 = (^({3{((2'd3))}}>>(&((~(a2?b3:b0))!=(b3<=b4)))));
  assign y13 = (~&(3'd6));
  assign y14 = {2{{(^{3{a0}}),(|(~&{b5,a4,a1}))}}};
  assign y15 = (5'd5);
  assign y16 = (+({3{b0}}>={{2{b0}},(+p0)}));
  assign y17 = (~^a4);
endmodule
