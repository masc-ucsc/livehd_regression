module expression_00360(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'sd2)<<<(-5'sd1))!=((3'sd1)-(-2'sd0)));
  localparam [4:0] p1 = {4{{1{((-5'sd14)>>>(5'd13))}}}};
  localparam [5:0] p2 = ((~|(~^(3'd1)))*((3'd3)<=(-2'sd0)));
  localparam signed [3:0] p3 = (((4'd4)-(2'd0))||{(3'd1),(2'd3),(-4'sd6)});
  localparam signed [4:0] p4 = {((3'd4)&(|(2'd2)))};
  localparam signed [5:0] p5 = (4'd11);
  localparam [3:0] p6 = (2'd1);
  localparam [4:0] p7 = {1{(^{((2'd3)<=(5'd2))})}};
  localparam [5:0] p8 = ({4{(4'd4)}}||{3{(3'sd2)}});
  localparam signed [3:0] p9 = {1{{1{(4'd8)}}}};
  localparam signed [4:0] p10 = ((!(6'd2 * (3'd2)))?(~^(((5'sd2)?(2'd1):(3'sd2))>=(~&(2'd0)))):(((4'sd4)>=(-2'sd0))?(5'd17):((5'sd8)||(-3'sd0))));
  localparam signed [5:0] p11 = (^(5'd21));
  localparam [3:0] p12 = {3{((2'd1)<(-4'sd5))}};
  localparam [4:0] p13 = ({(5'sd8),(2'd1)}||((5'sd1)^~(2'd0)));
  localparam [5:0] p14 = (!(((3'd7)?(-3'sd2):(3'd0))?(~&(-{(2'd3)})):((2'd3)?(4'sd2):(4'd12))));
  localparam signed [3:0] p15 = {{(3'd3),(2'd3)},((3'd7)>(5'sd8))};
  localparam signed [4:0] p16 = ((~^(!(&(((-5'sd11)>(4'sd0))!==(~&(5'sd9))))))>>>(-5'sd10));
  localparam signed [5:0] p17 = ((5'sd12)&&(3'd3));

  assign y0 = (+(~^$signed((-3'sd1))));
  assign y1 = {3{({4{b4}})}};
  assign y2 = {(a4==a5),(p1>b2),(b3>>>a5)};
  assign y3 = ((b3^b0)|(a0>=a0));
  assign y4 = (4'd7);
  assign y5 = (((b3)!={a1})>>{(a1||a5),(-a1)});
  assign y6 = ((2'd0)&({b2,a2}|(4'd7)));
  assign y7 = (({2{p5}}<<(2'd2)));
  assign y8 = {4{$signed((5'd27))}};
  assign y9 = {2{(5'd3)}};
  assign y10 = (&(((a2^~b3)!=(~|(p17||b0)))||{{b0,p16,a0},(b0+b5)}));
  assign y11 = (((p17&&p16)^~(a1&p15))-((p2<<b5)||(a5|p7)));
  assign y12 = (-2'sd1);
  assign y13 = (((4'd2 * (a2?b2:a1))==={3{a4}})>=(((p16?a5:a5)>>(b1?p14:a2))+(a3?a3:b3)));
  assign y14 = ({1{(3'd7)}}!==((a3!=a4)?{3{b3}}:(a4>>>a0)));
  assign y15 = ({3{(-2'sd0)}}!==((3'sd0)?(a0?a4:a4):(5'sd8)));
  assign y16 = (~&((a5?a4:a3)?(b0):(a0)));
  assign y17 = $unsigned((4'd2 * (-(&p8))));
endmodule
