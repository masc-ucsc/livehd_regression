module expression_00799(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^({(+(~(-3'sd3))),(~{(2'd2)})}|{((4'd9)||(3'd0)),((-3'sd3)==(-3'sd1)),((5'd3)<=(5'd10))}));
  localparam [4:0] p1 = {((~^((2'sd0)^~(5'd4)))+(&(|(&(3'd5))))),(+(((5'sd8)&(3'sd0))>(+(^(5'd10)))))};
  localparam [5:0] p2 = (((2'd2)?(5'd20):{(5'd16),(-5'sd12),(3'd1)})?{3{((-2'sd0)?(-2'sd1):(5'sd8))}}:{((-5'sd14)?(4'sd3):(3'd6))});
  localparam signed [3:0] p3 = {(~^({((3'd0)>(5'd5)),(~|(4'sd5)),((-3'sd3)?(3'd4):(5'sd13))}?((~(5'd24))?(+(5'd14)):(4'sd4)):(((2'd3)?(2'd0):(5'd6))===((-2'sd0)<(2'd2)))))};
  localparam signed [4:0] p4 = (4'd15);
  localparam signed [5:0] p5 = (((-4'sd7)||(-2'sd1))%(4'd4));
  localparam [3:0] p6 = (((-5'sd11)==(3'd7))+(5'd9));
  localparam [4:0] p7 = (((2'd1)?(5'sd2):(4'sd4))?((5'd14)<(5'd1)):(&(3'd3)));
  localparam [5:0] p8 = (+(~^(~(((~^(3'd1))<(+(5'd27)))+{3{(~|(2'sd0))}}))));
  localparam signed [3:0] p9 = (5'sd13);
  localparam signed [4:0] p10 = {(4'd0)};
  localparam signed [5:0] p11 = (+{({(3'd4)}==((3'sd2)<=(-5'sd3))),({(-5'sd3)}-{3{(5'sd7)}})});
  localparam [3:0] p12 = (((3'd6)>(4'd9))&(^(2'd0)));
  localparam [4:0] p13 = {4{(3'd4)}};
  localparam [5:0] p14 = (((~(5'd19))?((2'd2)^(5'd3)):((3'd0)?(3'sd1):(5'd3)))>=(!(~&((-(2'd3))&((4'sd5)|(3'd3))))));
  localparam signed [3:0] p15 = (~&(~&(|(^(-5'sd7)))));
  localparam signed [4:0] p16 = (~|(~|(((3'sd1)+(3'd0))%(4'sd2))));
  localparam signed [5:0] p17 = ((((-3'sd3)%(2'sd1))?((5'sd14)?(5'd16):(-4'sd6)):((2'sd1)>>(2'd3)))>(((-4'sd5)?(2'sd0):(3'd1))?((3'sd3)?(-3'sd2):(3'sd1)):((-3'sd1)-(4'd1))));

  assign y0 = {(~{((b4<<b1)!==(a4!=b5)),((b1>>b3)==(p13==a1)),{({b3,a3}>>>{a0})}})};
  assign y1 = (5'd22);
  assign y2 = {a2,b5};
  assign y3 = {4{$signed((p14>>p8))}};
  assign y4 = (!({1{{(&((2'd2)?$unsigned({a2,p8,b5}):{(2'd0),(+a1),(3'd6)}))}}}));
  assign y5 = (2'sd0);
  assign y6 = (({{(p2?p10:p14)},(p17?p9:p8)})<{{4{p12}},{p2,p2,p9},{2{p13}}});
  assign y7 = ((|$signed($unsigned(((a0<b2)!=(p9>>>p11))))));
  assign y8 = ({2{{1{(5'd10)}}}}!==($signed((-4'sd5))^(b5<b1)));
  assign y9 = (5'd2 * (^(p13>=p8)));
  assign y10 = ((~|b4)/a3);
  assign y11 = {({a4,p13,a2}?(b1?b2:a5):(~|{a1,b3}))};
  assign y12 = {{({{2{(p8?p15:p3)}}}?(!((p3?p3:p13))):(~^{{1{p14}},(p5?p6:p16),$unsigned(p5)}))}};
  assign y13 = {(|{{(~&(^(&(5'd24))))},(&(-(^(~(~|p11))))),(&{(~^(^(~|p7)))})})};
  assign y14 = $unsigned((-(((~^$unsigned(((~|$signed(p6))>(a4===a5)))))-$signed($signed(((-(b4===b2))&&$signed($signed(p15))))))));
  assign y15 = ($unsigned((+(^p3)))||((-p1)^$signed(b2)));
  assign y16 = {{{(|{p5,b5})}},{((^b1)|{p1,p10})},({p15,p0}<=(a4!==a5))};
  assign y17 = {{(^((~^(5'd25))?{p4,a1}:$signed((p0&p13))))},(^$signed((4'sd7)))};
endmodule
