module expression_00289(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((4'd7)^(5'd29)),{(4'd5),(3'sd0),(4'sd1)},(&{(5'sd12)})};
  localparam [4:0] p1 = ({3{(5'd3)}}?((3'sd1)||(2'sd1)):((-3'sd0)?(5'sd1):(3'd6)));
  localparam [5:0] p2 = {1{((-5'sd4)?(3'd2):(4'd2))}};
  localparam signed [3:0] p3 = (2'd2);
  localparam signed [4:0] p4 = ({3{(3'd4)}}?((2'd0)+(5'd24)):{1{{2{(2'd1)}}}});
  localparam signed [5:0] p5 = ((+((-3'sd0)&(2'sd0)))<=((3'd6)<=(-3'sd3)));
  localparam [3:0] p6 = ((2'd2)*(4'sd3));
  localparam [4:0] p7 = (5'sd8);
  localparam [5:0] p8 = {({4{(4'd10)}}|((3'd5)<<(3'sd1))),{1{({4{(3'd5)}}&&((-3'sd2)&(4'd7)))}}};
  localparam signed [3:0] p9 = (^(~|(3'sd1)));
  localparam signed [4:0] p10 = (((-4'sd5)^((3'd7)?(4'd0):(-4'sd6)))?{((4'd15)^~(-2'sd0)),((2'sd1)!=(-4'sd2))}:(2'd0));
  localparam signed [5:0] p11 = (((4'd14)?(-2'sd0):(5'd6))?((-4'sd1)===(2'sd0)):(-2'sd0));
  localparam [3:0] p12 = ({1{(~(2'sd1))}}?{3{(3'd3)}}:((3'd3)^(-4'sd0)));
  localparam [4:0] p13 = (((+(-4'sd4))?((3'd7)|(2'd0)):(-3'sd1))>=(+(|(~((-3'sd3)?(2'd0):(3'sd3))))));
  localparam [5:0] p14 = {1{(-5'sd6)}};
  localparam signed [3:0] p15 = {(4'd8),((-2'sd0)<=(4'd2))};
  localparam signed [4:0] p16 = ((-3'sd1)?(-4'sd6):(3'd2));
  localparam signed [5:0] p17 = {(-4'sd0)};

  assign y0 = ((!$signed((-2'sd1)))?((~(p14||p10))>>(4'd2 * p2)):$unsigned((~(p1?p3:p17))));
  assign y1 = ({4{{p1,b1,b3}}}<<<$signed($unsigned($unsigned((-$signed(((b3||p10))))))));
  assign y2 = ($signed($signed($signed((2'd0))))^({p11,a4,p13}<<<((5'd28)|(p9>p4))));
  assign y3 = (~&(~|(+(~(!(^(-(~|(+(!(~|p3)))))))))));
  assign y4 = {3{{4{p14}}}};
  assign y5 = (({1{{{{p7,p5},$unsigned(p16)}}}})+{{p8,p5,p2},$signed({p4,p10})});
  assign y6 = (5'sd10);
  assign y7 = ({2{({a4,b0,a2}?(~b5):(~&a3))}}-{3{(p3&&b5)}});
  assign y8 = (3'd5);
  assign y9 = (b2?a2:a3);
  assign y10 = {3{(b4?a3:a1)}};
  assign y11 = (+(|(p14<<<a2)));
  assign y12 = {4{(!p17)}};
  assign y13 = {1{(((p16<=p1)?{3{p17}}:{3{a3}})?{{2{b5}},(p7?p14:p1),(a4&&p12)}:{3{{1{b2}}}})}};
  assign y14 = (5'd2 * (b1!==b1));
  assign y15 = ($unsigned(a1)%a3);
  assign y16 = ((4'sd3)<{2{b3}});
  assign y17 = {3{(-4'sd3)}};
endmodule
