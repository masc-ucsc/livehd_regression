module expression_00522(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+(((5'd27)|(3'd5))||((5'sd9)>>(3'd1))))===((~|(5'd5))^(^(-5'sd9))));
  localparam [4:0] p1 = (((-3'sd2)?(2'd0):(3'sd1))>((6'd2 * (2'd2))&(&(3'sd3))));
  localparam [5:0] p2 = (-(2'sd0));
  localparam signed [3:0] p3 = {(2'd3),(4'd8),(-4'sd4)};
  localparam signed [4:0] p4 = ((+(((5'd12)==(5'd30))&((2'd3)?(5'd28):(4'sd2))))||((~^(4'sd2))===((2'd1)>(2'sd1))));
  localparam signed [5:0] p5 = {(|({2{(4'sd6)}}|((-5'sd9)===(3'd6)))),({2{(2'd2)}}==((5'sd0)>=(4'd15)))};
  localparam [3:0] p6 = (5'sd1);
  localparam [4:0] p7 = (-4'sd6);
  localparam [5:0] p8 = (5'd16);
  localparam signed [3:0] p9 = ({(-5'sd7),(3'sd2),(4'sd0)}!=({(3'd3)}<<{2{(3'sd0)}}));
  localparam signed [4:0] p10 = ((((~&(3'sd2))<=(~|(-2'sd1)))<<({4{(-3'sd3)}}<<(~&(2'd3))))>>({4{(3'sd2)}}^~{2{((5'd15)!=(2'd3))}}));
  localparam signed [5:0] p11 = (+{3{(2'd3)}});
  localparam [3:0] p12 = ({3{(4'd14)}}<(~^(-5'sd4)));
  localparam [4:0] p13 = ({(4'd15),(-4'sd3)}=={(4'd12),(4'd4)});
  localparam [5:0] p14 = ({(3'sd1),(3'sd0)}?((-2'sd0)+(5'd10)):{(-4'sd2),(3'd3)});
  localparam signed [3:0] p15 = (4'd2 * {1{(|(4'd8))}});
  localparam signed [4:0] p16 = (((-3'sd1)?(-4'sd1):(-4'sd7))?((2'd2)?(3'sd1):(3'd2)):(~|(^(-2'sd0))));
  localparam signed [5:0] p17 = ((-4'sd3)<<<((3'sd0)?(2'd1):(2'sd0)));

  assign y0 = (5'd15);
  assign y1 = ((!{{1{a1}}})<{a4,a2,p9});
  assign y2 = (3'd0);
  assign y3 = ((~&(!((^p10)?(~|p14):(-4'sd0))))^~((&p15)?(4'sd1):(|p6)));
  assign y4 = $unsigned(($unsigned(b4)%a3));
  assign y5 = (({a5,p6,p0}<<(5'd2 * (-a2)))<<((~(a1!=a3))==={(b5>>a1)}));
  assign y6 = ({4{(a0)}}^~(((b1-b0)==(|b5))+$unsigned({a3,b4,p5})));
  assign y7 = (b0?b4:a0);
  assign y8 = (4'd3);
  assign y9 = (3'd1);
  assign y10 = {3{(p9)}};
  assign y11 = ((p15^p11)&&(p10));
  assign y12 = (((p1<<p4)>(b0>>>b3))+{{p9,b3,p15},(b1!==a3),(b0!==a5)});
  assign y13 = {4{$unsigned(p8)}};
  assign y14 = (~^({1{$signed(({1{p12}}>={1{p3}}))}}&{3{{2{p8}}}}));
  assign y15 = (p1<<<p4);
  assign y16 = (~{3{{1{(p1>=p4)}}}});
  assign y17 = $signed((2'd3));
endmodule
