module expression_00497(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^{(&(~^{(4'sd0),(-2'sd1),(4'd11)})),(~&((4'sd3)?(3'd5):(2'd1))),(~^(^((-3'sd2)?(4'd6):(2'd0))))});
  localparam [4:0] p1 = (((-2'sd0)*(4'sd5))/(5'd14));
  localparam [5:0] p2 = (&({(5'd29)}!=(5'd2 * (2'd0))));
  localparam signed [3:0] p3 = (((2'sd1)<<(5'd25))*((2'sd1)<(-2'sd0)));
  localparam signed [4:0] p4 = {2{(!(+({2{(2'd2)}}>>(~&((5'd0)<=(4'd12))))))}};
  localparam signed [5:0] p5 = (((-5'sd15)^~(4'sd5))&&((4'd13)+(2'd3)));
  localparam [3:0] p6 = ((-5'sd0)?(5'd1):(5'd26));
  localparam [4:0] p7 = ({1{(4'd3)}}==(((3'sd2)>>((5'd14)!=(2'd3)))!==(-((2'd0)<(4'sd0)))));
  localparam [5:0] p8 = {(&(3'sd2))};
  localparam signed [3:0] p9 = (((-2'sd0)>>>(5'sd3))*(+(-2'sd0)));
  localparam signed [4:0] p10 = {((3'd7)&&(3'd0)),(|((4'sd3)^~(4'sd5))),((3'sd2)>(2'sd0))};
  localparam signed [5:0] p11 = (((-5'sd6)?(5'sd6):(2'd0))?(^((2'sd1)|(4'd1))):(+((2'sd1)+(3'd2))));
  localparam [3:0] p12 = {2{{1{(+((-3'sd2)?(-3'sd3):(5'd19)))}}}};
  localparam [4:0] p13 = ((4'd14)*((3'd2)!==(4'd12)));
  localparam [5:0] p14 = ((((4'd5)&(2'd3))>=(|((2'd3)!==(5'd12))))^(~^(&(~&((-5'sd5)%(-5'sd7))))));
  localparam signed [3:0] p15 = (+(((2'd2)?(4'd1):(4'd9))?(~((5'd21)>=(2'd1))):(-3'sd3)));
  localparam signed [4:0] p16 = {3{(-2'sd1)}};
  localparam signed [5:0] p17 = (5'sd5);

  assign y0 = ({4{a3}}>>{2{{p12}}});
  assign y1 = (a2<<p6);
  assign y2 = {2{(2'd3)}};
  assign y3 = (~&{(&(~|(-(+{(~&a2),{a3},(~&a5)})))),(-(~(5'd29)))});
  assign y4 = ({4{p1}}!={4{p1}});
  assign y5 = $signed((p13||a4));
  assign y6 = {2{((b5?p17:b2)?(a1?b3:p11):{2{p12}})}};
  assign y7 = ((^((~&$signed({b4}))===((a3>=a2)|(~&a0))))!=(~^(-4'sd1)));
  assign y8 = (~(5'd2 * (p14==p0)));
  assign y9 = (~&(^(!{1{{2{(&(~((&a3)==(~|b5))))}}}})));
  assign y10 = ((a4>=b1)<<(a3&a5));
  assign y11 = {(~&p12),(~&p11)};
  assign y12 = ({({p12,a2,b4}&&(a2===b2))}&&((~^(b3<<b0))!==(~^{b1,b2,a5})));
  assign y13 = ({2{(p14<=b4)}}?{2{(p1?p17:p0)}}:((p5?p2:a2)^(p17?b5:p8)));
  assign y14 = {((^(a5?b1:b1))),(+(6'd2 * {a2,a0,p12})),(-(&(^(!(~^a0)))))};
  assign y15 = {4{a4}};
  assign y16 = (~&$signed({4{{p15,p14}}}));
  assign y17 = {{{(p17^p3),(p15+p4),(p17^p7)}},{((a3&p0)>>>(p2>a5))}};
endmodule
