module expression_00232(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{((+(2'd3))>>>(!(2'sd0)))}}-(~^(~{2{{4{(3'd7)}}}})));
  localparam [4:0] p1 = (2'd3);
  localparam [5:0] p2 = (((3'd2)^(4'd0))^(!((-4'sd1)?(2'sd1):(2'd2))));
  localparam signed [3:0] p3 = (4'sd7);
  localparam signed [4:0] p4 = (5'd3);
  localparam signed [5:0] p5 = (2'd1);
  localparam [3:0] p6 = ((5'sd10)-(2'd0));
  localparam [4:0] p7 = {{4{{(5'd18)}}},{1{{{1{(4'd12)}},{(3'd6),(-5'sd6)},{(-4'sd0)}}}}};
  localparam [5:0] p8 = {{2{{3{(5'sd4)}}}}};
  localparam signed [3:0] p9 = {2{{(4'd15),(-2'sd0),(2'sd0)}}};
  localparam signed [4:0] p10 = (&(-(-3'sd2)));
  localparam signed [5:0] p11 = ((|((3'sd0)>>>(5'd31)))?((2'sd0)?(-3'sd1):(-3'sd2)):((|(3'sd1))<=((-4'sd4)?(-5'sd2):(4'd3))));
  localparam [3:0] p12 = ((2'd0)?(5'd31):(2'd3));
  localparam [4:0] p13 = (~(~&{((~&{(~^(-5'sd6)),(~&(4'sd3)),(~^(4'd2))})>>(-(-(-((4'd15)^~(3'd5))))))}));
  localparam [5:0] p14 = ((4'd11)>>(5'd31));
  localparam signed [3:0] p15 = ({1{((2'sd0)?(4'd15):(3'd4))}}?{1{(~|(&(2'd2)))}}:{1{((3'sd3)?(4'd6):(5'sd12))}});
  localparam signed [4:0] p16 = (~&{2{(3'd7)}});
  localparam signed [5:0] p17 = ((-3'sd2)||(2'sd1));

  assign y0 = (!(((a5%a4)?(^(a4?a2:a3)):(a3?a5:a3))&((~^(b4>a2))===(2'd0))));
  assign y1 = ((+(!{($unsigned($unsigned((2'd0)))!==((~^(~&{b4}))))})));
  assign y2 = (!({{2{a3}},(|{1{p0}}),{(~|p3)}}>>(|{4{{p7,b5}}})));
  assign y3 = (($unsigned(({a5,b0}<<<{p7,p8,b2}))-$signed({p17,b3,a5})));
  assign y4 = (5'sd15);
  assign y5 = (|{2{($unsigned({{b3},(~|p9)})>>>(-{(~&b0),{b5,p13}}))}});
  assign y6 = (((p17&a0)?(p12?b0:p9):(~|p2))?((b1>=a1)<(a3>b5)):{(b3?b4:b2),(p7?a1:p1),(a2!==b0)});
  assign y7 = ({4{a0}}||(&b3));
  assign y8 = ((-4'sd5));
  assign y9 = (~|(^((^((b0!=b2)<=(b3<<b4)))<=((b4/b0)&&(-(!a4))))));
  assign y10 = ((3'd6)<(+(~|$unsigned($unsigned((^(4'd2 * $unsigned(p1))))))));
  assign y11 = ({a5,a3,a4}^(p17>p9));
  assign y12 = (p11%p16);
  assign y13 = $signed($signed($signed($unsigned(({3{p14}})))));
  assign y14 = {3{p6}};
  assign y15 = (~^b4);
  assign y16 = {{((p13?p1:p15)?(-2'sd0):$signed(p16)),((p16)?{2{p6}}:(3'd4))}};
  assign y17 = (((p7>b3)?((b4^p8)):{{a3}})|(2'sd1));
endmodule
