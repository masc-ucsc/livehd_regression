module expression_00081(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd0)?{(4'd11),(2'd3)}:((4'd7)?(-2'sd0):(-3'sd0)));
  localparam [4:0] p1 = (((-5'sd13)>=(3'sd3))&&((-5'sd3)^~(4'sd1)));
  localparam [5:0] p2 = ((((-5'sd13)?(5'd14):(3'd1))?{(2'sd0),(-5'sd4),(-2'sd0)}:((2'sd0)>>(2'sd0)))===(((-3'sd0)^(3'd1))|((5'sd15)+(2'd1))));
  localparam signed [3:0] p3 = (~&(((3'd3)?(-5'sd12):(5'sd6))===(^((5'd10)?(3'd5):(3'd6)))));
  localparam signed [4:0] p4 = (4'd10);
  localparam signed [5:0] p5 = ({4{(2'sd0)}}<(+{4{(-4'sd0)}}));
  localparam [3:0] p6 = ((4'sd0)>=(-3'sd0));
  localparam [4:0] p7 = (!(!(!(!((4'sd1)+(-3'sd1))))));
  localparam [5:0] p8 = (((3'sd2)<=(2'd2))?((-3'sd0)>>>(4'sd6)):{3{(2'sd0)}});
  localparam signed [3:0] p9 = {(4'd13),(-2'sd1),(5'd17)};
  localparam signed [4:0] p10 = (((2'd1)?(3'd4):(4'd6))?(&((3'd4)?(3'd7):(5'd31))):((5'sd11)?(4'sd6):(4'd8)));
  localparam signed [5:0] p11 = (+{1{(~&(3'sd1))}});
  localparam [3:0] p12 = (((-4'sd7)?(5'd20):(3'd7))?((3'sd1)<(4'd2)):(&(-5'sd2)));
  localparam [4:0] p13 = {({(4'd14),(2'd2)}|{4{(4'd7)}}),{(-(3'd6)),((4'd0)?(-2'sd1):(2'd3))},(~({3{(3'd3)}}>={(3'd7),(5'd28),(5'd1)}))};
  localparam [5:0] p14 = (~|((-{3{(2'd0)}})^~(((3'sd1)==(2'd3))!={(4'sd2),(4'd10),(4'd1)})));
  localparam signed [3:0] p15 = (-5'sd9);
  localparam signed [4:0] p16 = (((-3'sd0)!=(2'd0))?((4'sd7)===(5'd17)):((-2'sd0)<<(5'sd15)));
  localparam signed [5:0] p17 = {{(((3'd2)?(3'd3):(2'sd0))>>>((-3'sd0)?(3'd1):(-3'sd3))),{((3'sd0)-(-3'sd1)),((2'd1)!=(3'sd2))},(((5'sd15)|(4'sd0))<={(4'sd0),(5'sd14),(2'd0)})}};

  assign y0 = (((p14&&p5)&(5'd2 * p14))=={4{p14}});
  assign y1 = (({(b1>p14)}>{p17,a5,b4})|(6'd2 * {(~|p8)}));
  assign y2 = (~|(|(!(|(!(!(~|(&(~(&(~(|(&(+(-a4)))))))))))))));
  assign y3 = ((&b2)<=(+p4));
  assign y4 = (+(((a2^p5)==(b5>p5))>=({p8,p16}!=(5'd26))));
  assign y5 = ({2{b5}}?$signed(b1):(a1<<a4));
  assign y6 = (4'd0);
  assign y7 = $signed((4'sd3));
  assign y8 = ((p0?a3:a0)?(p8&&b0):$unsigned((5'd13)));
  assign y9 = ((|$unsigned({b4,a2,a4}))?{{p13,a0,p8},(3'sd2),{b0,p6,p11}}:(~$signed((-(b4?a2:p7)))));
  assign y10 = {3{{p7,a3}}};
  assign y11 = {a0,p8,a5};
  assign y12 = (((p2<b1)&&(p14==p3))+((p15%p5)^~(p16|b2)));
  assign y13 = $signed((~^(~(2'd3))));
  assign y14 = ({4{p5}}>>>{(p13+p4)});
  assign y15 = (&p9);
  assign y16 = ((~(4'd14))?(|((p5?p9:b3))):(b0?p5:p16));
  assign y17 = ((b5!=p4)^~{2{a4}});
endmodule
