module expression_00042(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({(2'd0)}<=((-4'sd0)>>(3'd3)))===({(4'sd6),(4'd1)}<((2'd1)+(-4'sd3))));
  localparam [4:0] p1 = (~&((&(|(^(2'd0))))<<<(5'd31)));
  localparam [5:0] p2 = {((3'd1)==(4'd2))};
  localparam signed [3:0] p3 = (&(+(5'd27)));
  localparam signed [4:0] p4 = (5'd7);
  localparam signed [5:0] p5 = (((2'sd1)^(3'd3))===((-4'sd3)^(4'sd5)));
  localparam [3:0] p6 = {3{(((4'd11)?(-5'sd0):(2'd1))?((2'd3)!=(-5'sd6)):(!(-2'sd1)))}};
  localparam [4:0] p7 = (4'sd0);
  localparam [5:0] p8 = {((~^(2'd3))>=(~^(3'sd0))),(~&{(~|(-4'sd6))}),{{(5'd8),(2'sd1),(2'd0)}}};
  localparam signed [3:0] p9 = (({2{(2'd3)}}?(~&(4'sd4)):{1{(-5'sd1)}})?{2{{3{(-3'sd3)}}}}:{2{{4{(-4'sd5)}}}});
  localparam signed [4:0] p10 = (~^((4'sd6)?(-4'sd1):(2'sd0)));
  localparam signed [5:0] p11 = (5'd1);
  localparam [3:0] p12 = ((((-5'sd12)==(4'd2))^~((3'sd3)&(5'd30)))?((5'sd11)?(4'sd7):(4'd7)):((-2'sd0)?(2'sd1):(-4'sd6)));
  localparam [4:0] p13 = {{(3'sd1),(2'd3)},{(4'd13),(4'd5),(-2'sd0)}};
  localparam [5:0] p14 = {3{{{(5'sd0),(3'd0)},{(5'sd15),(3'd7),(5'd1)}}}};
  localparam signed [3:0] p15 = (({(5'sd8),(4'd2),(-4'sd3)}^((4'sd4)<<<(-2'sd1)))>>>{2{((4'd3)&&(2'sd1))}});
  localparam signed [4:0] p16 = (5'd21);
  localparam signed [5:0] p17 = {(4'sd7),{{(4'd6),(5'd15)},((-2'sd0)&(5'd21))},(4'd10)};

  assign y0 = (+((~&(p12!=p3))&((|p11)<=(5'd2 * p2))));
  assign y1 = (~(+((-3'sd3)*(b0-p2))));
  assign y2 = (-3'sd0);
  assign y3 = (((5'd26)/p0)>>>((3'd5)>>>((b0?a3:a5)!==(a3&b4))));
  assign y4 = (&(a5>>>b0));
  assign y5 = (~{3{{1{{4{a2}}}}}});
  assign y6 = (5'd0);
  assign y7 = (((a3-p4)?(a5|b0):(5'sd13))?((-2'sd1)>(p10?p2:a5)):((2'd3)?(a0!==a5):(a1/p4)));
  assign y8 = $signed((!{(~|((b0?a4:p14)?$unsigned(a0):(a0^~b4)))}));
  assign y9 = ((|(b5!=a0))===((~|a0)>>>(^a2)));
  assign y10 = (((~&{3{a2}})<(p9^~p11))!=({2{p17}}&&(a2||p11)));
  assign y11 = {p11,b3};
  assign y12 = ((6'd2 * (~&(&b0)))>>>(~^((b0!==a4)<<<(b1))));
  assign y13 = (a0||p6);
  assign y14 = (({p6,b2,p17}?(a5===b3):(p3<<b1))-((~^{a5})^(a5!==a0)));
  assign y15 = (~&(-$unsigned((b0>=b0))));
  assign y16 = {4{p10}};
  assign y17 = {1{{1{p4}}}};
endmodule
