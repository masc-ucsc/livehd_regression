module expression_00688(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(!(~|({2{((2'sd1)===(4'd13))}}==={2{(-(3'd0))}}))));
  localparam [4:0] p1 = {1{(!(~&{(~(!{2{(2'd0)}})),{{2{(-5'sd11)}},{(-2'sd0),(4'sd7),(3'd1)}},{(3'd6),(5'sd11),(4'd13)}}))}};
  localparam [5:0] p2 = {1{{1{(-4'sd6)}}}};
  localparam signed [3:0] p3 = ((4'sd0)?(3'd4):(-3'sd2));
  localparam signed [4:0] p4 = {4{((4'sd1)||(2'd3))}};
  localparam signed [5:0] p5 = (&{3{((~|(4'd6))!=={4{(2'sd1)}})}});
  localparam [3:0] p6 = (-3'sd2);
  localparam [4:0] p7 = ({(~|(4'd7)),{(4'd11)},{(2'd1),(5'd4)}}?({1{(-5'sd0)}}>((-5'sd8)>(5'd24))):{(-(2'd3)),((-2'sd1)<<<(-2'sd1))});
  localparam [5:0] p8 = {2{(+(((5'd16)-(3'd4))|((3'sd1)>(2'd3))))}};
  localparam signed [3:0] p9 = {3{{2{(3'd6)}}}};
  localparam signed [4:0] p10 = {3{((-2'sd0)<=(-4'sd1))}};
  localparam signed [5:0] p11 = ((2'd1)?(5'd7):(2'sd1));
  localparam [3:0] p12 = ((^(5'd17))?((2'd2)>=(2'd1)):((3'd6)<=(4'd4)));
  localparam [4:0] p13 = ((((-3'sd1)>>(2'sd1))&&((-4'sd1)&&(5'd30)))!==({1{(~|(2'sd1))}}>=((2'sd0)!==(2'd0))));
  localparam [5:0] p14 = ((2'd2)||(4'sd6));
  localparam signed [3:0] p15 = ({(4'sd0)}?((2'd1)?(3'sd0):(2'd3)):{1{(4'sd2)}});
  localparam signed [4:0] p16 = (((-5'sd9)-(2'sd1))?((-5'sd5)!==(4'sd4)):((4'd6)>=(4'd4)));
  localparam signed [5:0] p17 = (((2'd0)?(-3'sd2):(4'd11))<<<(^(3'd4)));

  assign y0 = ({(+{p16,a0}),((+a3)),(-(p4))});
  assign y1 = (((a5==b4)>>>(p10+a4))>((a1!==a0)^(b3==a1)));
  assign y2 = (^(-(-4'sd0)));
  assign y3 = (!((3'sd3)));
  assign y4 = ((!(p3?p7:p14))?(3'd6):{2{p4}});
  assign y5 = ((-2'sd1)&(5'd2 * (p1<<<p8)));
  assign y6 = (5'd24);
  assign y7 = $signed($signed(($signed((a1?p16:p2))<<{{p15},(p8!=p10)})));
  assign y8 = ((5'd28)||(!(3'd0)));
  assign y9 = ((^((&(p6?p3:p0))))||(-4'sd6));
  assign y10 = ((p16|p11)*$unsigned((a5+p8)));
  assign y11 = (((p6?b4:b4)?$signed($unsigned(a2)):(a4?b4:a3)));
  assign y12 = (2'sd0);
  assign y13 = ({a3,a3,b4}>={b0,a4});
  assign y14 = (~|(((~|(a1^a5))^(2'd0))&(5'd2 * (b1^p0))));
  assign y15 = {2{{{3{b3}},{4{a2}},{4{b1}}}}};
  assign y16 = (+(3'd7));
  assign y17 = $unsigned({3{$signed(a2)}});
endmodule
