module expression_00708(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(3'd0));
  localparam [4:0] p1 = (~^((3'd5)?(3'sd0):(4'sd0)));
  localparam [5:0] p2 = (~|{(-3'sd1)});
  localparam signed [3:0] p3 = (~^(|{2{(-5'sd8)}}));
  localparam signed [4:0] p4 = {2{{((-2'sd1)===(3'd0)),{(2'd1),(2'd0)},(6'd2 * (4'd14))}}};
  localparam signed [5:0] p5 = (3'd3);
  localparam [3:0] p6 = ({{1{(+(3'd0))}},{3{(2'sd0)}}}||({4{(-4'sd7)}}&(|((3'd1)>>(5'd19)))));
  localparam [4:0] p7 = (((4'sd5)?(5'd31):(5'd16))?{1{{2{(2'd2)}}}}:{3{(4'd14)}});
  localparam [5:0] p8 = (^(~|((|(2'sd1))?{(2'd2)}:(!(5'd15)))));
  localparam signed [3:0] p9 = ((2'sd0)*((4'sd2)!==(3'sd1)));
  localparam signed [4:0] p10 = ((|{4{(2'sd0)}})+(~&(3'd3)));
  localparam signed [5:0] p11 = ((5'd30)||(4'sd6));
  localparam [3:0] p12 = (4'd10);
  localparam [4:0] p13 = {{(((-2'sd0)&(5'd6))||((3'd2)<<<(-2'sd1)))},({(3'sd1),(3'sd0)}?((3'sd1)^(4'sd2)):(&(3'sd1)))};
  localparam [5:0] p14 = {(((!(-2'sd0))==((2'd2)?(5'd18):(4'sd7)))<<{3{((2'sd0)+(3'd5))}})};
  localparam signed [3:0] p15 = (&({(^(4'sd7))}?((2'd1)?(4'd13):(2'd0)):(~^(!(4'd5)))));
  localparam signed [4:0] p16 = ((5'd2 * {(3'd0),(2'd3),(3'd6)})||({(3'd0),(5'd29),(4'd4)}?((-2'sd0)==(-5'sd8)):(+(5'd14))));
  localparam signed [5:0] p17 = (~&((!{1{(!(5'sd14))}})==(~|(+((3'd4)<<(-5'sd13))))));

  assign y0 = {((^{b3,b1,b4})?{a5,a2,b2}:{(+b2)})};
  assign y1 = (b5?p14:a5);
  assign y2 = (b3!=a1);
  assign y3 = ((~&(p13?a2:p5))?$unsigned($unsigned(a0)):(-(p10?p3:a1)));
  assign y4 = ((((b3===a4)<=(p8>>>p3))==(5'd2 * (p0>>>b1)))<(((p14>p15)*(a3==p3))<<<((p6<=a4)/p16)));
  assign y5 = (((4'sd5)^(a4?p1:b4))?(3'd6):(3'sd0));
  assign y6 = (~^$signed((4'sd5)));
  assign y7 = ((a1?a2:b0)?{1{(b3?a5:b2)}}:(~(~^{2{a4}})));
  assign y8 = (((p9?p2:b2)<(p16?p4:p13))>>>((p8&p9)?(p3%p14):(p3==p14)));
  assign y9 = (+(^(|(~|(~^(b0<p5))))));
  assign y10 = {{{3{{4{p15}}}},{1{{4{b1}}}},{1{(&(!{p11,b3}))}}}};
  assign y11 = $signed({4{({1{b2}}<=(a3))}});
  assign y12 = {2{$signed(((+{1{(+$signed((&p13)))}})))}};
  assign y13 = (p5?b2:a1);
  assign y14 = $signed(({p15,b2}|{$unsigned(p2)}));
  assign y15 = {(|{4{p12}}),{(p6&&p0),{p5,p0,p1}},{{(p0||p13),(|p13),(~^a4)}}};
  assign y16 = (!($unsigned((p3+p4))&&(p15<=p1)));
  assign y17 = (p10?p16:p4);
endmodule
