module expression_00001(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'd7);
  localparam [4:0] p1 = ((-5'sd14)<(5'd1));
  localparam [5:0] p2 = ((-4'sd2)>>>(^(4'd0)));
  localparam signed [3:0] p3 = ((~^(3'd3))-(|{(4'd9),(5'd24)}));
  localparam signed [4:0] p4 = {2{((2'd3)>=(4'sd3))}};
  localparam signed [5:0] p5 = (({(3'd5)}^~((5'd30)+(3'd7)))<(((3'd7)<(4'd14))>=((-3'sd2)==(4'd15))));
  localparam [3:0] p6 = ((4'd1)?(2'sd0):(2'd3));
  localparam [4:0] p7 = (&{4{(-3'sd2)}});
  localparam [5:0] p8 = ({4{(2'd1)}}>>{3{(5'd13)}});
  localparam signed [3:0] p9 = (4'sd5);
  localparam signed [4:0] p10 = ((3'd4)===(((4'd2)===(5'd10))>(-3'sd3)));
  localparam signed [5:0] p11 = (((2'd0)?(3'd7):(2'sd0))?(2'sd1):((5'd8)?(5'd17):(5'd25)));
  localparam [3:0] p12 = (5'd0);
  localparam [4:0] p13 = (4'd2 * (3'd1));
  localparam [5:0] p14 = (((~^(2'd0))*((5'sd2)?(3'sd0):(5'd11)))|(|(|((4'd2)?(4'sd4):(2'd2)))));
  localparam signed [3:0] p15 = ((4'd2 * (+((3'd7)<<(3'd1))))===(((3'd7)&(-3'sd1))||((-5'sd6)*(2'd1))));
  localparam signed [4:0] p16 = (-(-(3'd5)));
  localparam signed [5:0] p17 = (~({(~^((2'sd0)>>>(-3'sd2)))}?{(5'd14),(5'sd9),(3'd0)}:(((2'd3)^(4'd5))!=(~|(3'sd0)))));

  assign y0 = (((&a1)^~(!a0))>>((-a5)>(^b1)));
  assign y1 = {((~^(|(b3<=p4)))&{(~^a0),(b3>a4)}),(-3'sd3)};
  assign y2 = {{(&(~a0)),{a5,p3,b5},(~^(~^p1))},(-$unsigned((~|$signed({(|b5),(!a1),(~^a4)}))))};
  assign y3 = (^((6'd2 * (~^$unsigned(b5)))|(+(!{2{{4{b0}}}}))));
  assign y4 = (p13<<<p10);
  assign y5 = ((^((~^p9)^{4{a5}}))?{3{(-2'sd0)}}:((~&(p5<=b2))>(3'sd0)));
  assign y6 = (~|(3'd3));
  assign y7 = (~(((a2-b1)%b4)<=((a0?b4:a3)>>>(b0?a3:a3))));
  assign y8 = ((~|(a3?p6:p5))?{a2,p13,a1}:(a4?p10:a1));
  assign y9 = ({4{(a5?a1:a2)}}?((a2||b1)?(b1-b3):{3{b0}}):((a2<=b4)===(a5?a3:a1)));
  assign y10 = (5'd22);
  assign y11 = (+(~^((6'd2 * (~^(&a0))))));
  assign y12 = (|{(~&{2{{(|(!a0)),{(b3!==a2)}}}})});
  assign y13 = {2{((-5'sd6)?(-5'sd15):(b2<<a5))}};
  assign y14 = (4'd1);
  assign y15 = {{4{p2}},(~&(|{2{p16}})),(&((p6<p5)>>>{p9,p3}))};
  assign y16 = {{{b3},{2{a3}},(b4==a3)},{({2{b0}}),$unsigned({4{b4}})}};
  assign y17 = (((~&b0)>>>(p0?p13:b1))!=(p12?p17:a3));
endmodule
