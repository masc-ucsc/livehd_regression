module expression_00225(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({2{(!{4{(5'sd10)}})}}||(-({2{(2'd3)}}?((-5'sd10)<(3'sd1)):{2{(2'd0)}})));
  localparam [4:0] p1 = {3{((-5'sd14)^~(4'd9))}};
  localparam [5:0] p2 = (({2{(-4'sd0)}}!==((2'sd1)-(4'sd7)))<{3{(+(2'd0))}});
  localparam signed [3:0] p3 = (5'd21);
  localparam signed [4:0] p4 = {((-3'sd0)+(-2'sd1)),(-4'sd2),(!(-4'sd0))};
  localparam signed [5:0] p5 = (~{2{{1{(^(+((-3'sd2)+(5'sd12))))}}}});
  localparam [3:0] p6 = (-5'sd0);
  localparam [4:0] p7 = ((-2'sd0)===(~&(|(-4'sd7))));
  localparam [5:0] p8 = {{(2'd1),(2'd1),(-4'sd0)},((3'd2)?(-4'sd0):(4'sd6))};
  localparam signed [3:0] p9 = (((2'd3)>>(5'sd4))===((-4'sd7)?(4'd2):(-5'sd7)));
  localparam signed [4:0] p10 = ({3{(5'sd0)}}!=(-((5'd0)>>>(-2'sd1))));
  localparam signed [5:0] p11 = {2{(4'd2 * ((4'd8)-(5'd25)))}};
  localparam [3:0] p12 = (-(({(-2'sd0),(3'd6)}&&{(2'sd0)})==(~&((5'd0)<=(4'd9)))));
  localparam [4:0] p13 = {(-5'sd4),(4'd7)};
  localparam [5:0] p14 = (!{1{(+((4'sd2)===(3'd5)))}});
  localparam signed [3:0] p15 = ((4'd2 * (3'd0))!={1{(-2'sd1)}});
  localparam signed [4:0] p16 = {2{(3'd0)}};
  localparam signed [5:0] p17 = ((&(((5'd0)^(2'sd0))?(|(3'd2)):((-5'sd0)*(-2'sd0))))<=(((5'sd4)*(4'sd5))!=((4'd9)?(3'd5):(2'sd0))));

  assign y0 = {{(!{a5}),((p1))},{(b1>>p8),{p16},(p6^~p8)}};
  assign y1 = ((&(5'd2 * (^(a0!==b1))))^~((~&(a2==a4))>=(!(~(~p7)))));
  assign y2 = (p9?p11:p4);
  assign y3 = {a3,a5};
  assign y4 = (~(~^{(5'd2 * b0),(~^a0),{p17,p1}}));
  assign y5 = ((p10?p9:p4)<(+(p2>=p6)));
  assign y6 = {2{({p17,p2,p15}^{p8,a1,p0})}};
  assign y7 = ((~|p12)!=(~|b5));
  assign y8 = {2{(4'd11)}};
  assign y9 = ((~b0)<<<$unsigned(b1));
  assign y10 = (&(-2'sd1));
  assign y11 = ((~(5'd17))>>{{a4,p15,p17},{p4,p12}});
  assign y12 = (5'd2 * (5'd2 * a2));
  assign y13 = ((~^$unsigned((p2)))!=$unsigned($signed($signed(a3))));
  assign y14 = (3'd5);
  assign y15 = (((a3?a4:b5)?$unsigned((p10?p3:a1)):(a3?b4:p7)));
  assign y16 = (a3);
  assign y17 = (+{((&b1)?(b4>>>b1):(|a5)),{(~((-b3)^~{a3,b1,a5}))},((~b5)?{a4,b4,b0}:{b5,b0})});
endmodule
