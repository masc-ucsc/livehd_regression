module expression_00744(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(-5'sd13),{(2'd2),(2'd2),(5'd26)}},{{(3'sd1),(3'd1),(-2'sd0)},(-5'sd2),(5'd14)}};
  localparam [4:0] p1 = {2{((&(2'sd1))?{4{(4'd5)}}:(~|(4'd6)))}};
  localparam [5:0] p2 = (~&(5'sd0));
  localparam signed [3:0] p3 = (((5'd24)?(-2'sd0):(3'sd0))?((3'sd3)?(-2'sd0):(3'd4)):((2'sd0)<<<(3'd6)));
  localparam signed [4:0] p4 = (~^(5'd20));
  localparam signed [5:0] p5 = (-5'sd0);
  localparam [3:0] p6 = ({4{(4'd2)}}?(((-3'sd2)||(3'd6))!=((5'd7)==(3'd3))):({1{(4'sd4)}}==={1{(5'sd1)}}));
  localparam [4:0] p7 = (((3'd2)-(5'd14))||(3'd2));
  localparam [5:0] p8 = (((3'd6)!=(3'd1))%(2'sd0));
  localparam signed [3:0] p9 = (~&(-3'sd2));
  localparam signed [4:0] p10 = ((&(4'd13))>=((3'd3)^~(4'd6)));
  localparam signed [5:0] p11 = (^((-{{(2'd1),(3'd7)}})?((5'd9)<<<(4'd9)):((5'sd6)?(5'sd7):(5'd1))));
  localparam [3:0] p12 = (5'sd15);
  localparam [4:0] p13 = (!(~((((4'sd7)==(-5'sd3))&&((5'd31)<=(4'd5)))!={1{(^((2'd2)!=(5'sd2)))}})));
  localparam [5:0] p14 = {1{({2{{((2'd1)||(2'd1))}}}<{2{((4'd8)&&(4'sd2))}})}};
  localparam signed [3:0] p15 = ((2'd1)?(((3'sd2)?(-4'sd1):(4'd11))>>>((4'sd3)?(-3'sd0):(5'd29))):(((3'sd2)?(-5'sd6):(-4'sd3))^~((4'd8)<=(2'd3))));
  localparam signed [4:0] p16 = (~{(2'd1),(5'd2 * {(3'd2),(3'd4),(4'd1)}),(|((2'd3)&(4'd10)))});
  localparam signed [5:0] p17 = ((((2'd3)>>(5'sd3))===(-2'sd1))&((-4'sd2)!=((4'sd6)>>(2'sd0))));

  assign y0 = (((a0^b5)));
  assign y1 = {(-5'sd14),{a5,b4,a4}};
  assign y2 = ($signed(p0)&&$unsigned(p3));
  assign y3 = (((2'd3)>(a4===a3))-(-4'sd4));
  assign y4 = (!$signed(p2));
  assign y5 = (((&b0)?(^b2):(a2))^~(-2'sd1));
  assign y6 = {3{((|a2)?(a0?b4:a0):(-b2))}};
  assign y7 = (&(((p3?p13:a2)|(p2==p7))?{(a1?p16:b2)}:((-b1)>>(a3?a0:b5))));
  assign y8 = ({(~b4),{b5,a1,a4}}!==(~|(5'sd5)));
  assign y9 = ((~^({a3,b1}==={b0,b4,a2}))>>>((a2^b5)>>{p16}));
  assign y10 = {3{(p6?p14:p1)}};
  assign y11 = (((3'd5))!==(-4'sd7));
  assign y12 = ((~p4)*$signed(a2));
  assign y13 = {((b4?a4:p3)?(a3<b3):{2{b2}}),{(-(a1||p12)),$signed((-4'sd7)),{4{a5}}}};
  assign y14 = (p17<<a0);
  assign y15 = {{(p7||p5),(~|(~&p4)),(p2?p0:p17)},(~&(3'd5))};
  assign y16 = (a2?b1:b1);
  assign y17 = (2'd2);
endmodule
