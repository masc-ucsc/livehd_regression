module expression_00272(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(+({1{(3'sd1)}}^((5'sd0)+(2'd1)))));
  localparam [4:0] p1 = (+(|{((~(+(5'sd12)))==={1{{(4'sd0)}}})}));
  localparam [5:0] p2 = (5'd31);
  localparam signed [3:0] p3 = (~&((((5'd28)||(-2'sd1))?((4'd10)&&(5'd14)):((4'd3)!==(2'sd0)))!==(((4'd10)==(-2'sd0))?((-4'sd4)<<(2'sd1)):(5'd2 * (4'd2)))));
  localparam signed [4:0] p4 = ((6'd2 * ((4'd15)>>(3'd6)))&&(((2'd2)<<(5'sd13))!=((5'sd10)===(2'd1))));
  localparam signed [5:0] p5 = ((((3'd5)==(5'd2))&((5'sd11)<=(-2'sd0)))=={((2'd2)?(3'd1):(3'sd3)),(2'd1),(3'd2)});
  localparam [3:0] p6 = (2'd3);
  localparam [4:0] p7 = (((2'd3)?(2'sd1):(5'sd12))?((5'sd11)?(3'sd3):(3'd5)):((4'd7)?(2'sd0):(5'sd8)));
  localparam [5:0] p8 = ((~((-4'sd0)===(-2'sd1)))-{4{(-4'sd3)}});
  localparam signed [3:0] p9 = ({4{(4'sd2)}}>{2{((3'sd1)==(4'd8))}});
  localparam signed [4:0] p10 = (~&(^((^(((3'sd3)?(3'd0):(3'd4))&(-(5'sd3))))&{1{{4{(5'd15)}}}})));
  localparam signed [5:0] p11 = {3{(-2'sd0)}};
  localparam [3:0] p12 = {3{((3'd6)<(4'd3))}};
  localparam [4:0] p13 = ((4'd10)>(5'sd4));
  localparam [5:0] p14 = {1{(-2'sd1)}};
  localparam signed [3:0] p15 = (3'd7);
  localparam signed [4:0] p16 = (3'sd3);
  localparam signed [5:0] p17 = {3{((5'sd14)?(4'd4):(3'd4))}};

  assign y0 = (~(~|(p10/p12)));
  assign y1 = {2{((5'sd0)?(b0!=b0):(2'sd1))}};
  assign y2 = (6'd2 * (~|{1{p8}}));
  assign y3 = (^$unsigned((&(&(!(~|((~^((~|p9)>=(|a1)))==(+(-(+(|(|b4))))))))))));
  assign y4 = (~|(a5!==b1));
  assign y5 = $signed((b0!==a3));
  assign y6 = {(!b1),(~^p11)};
  assign y7 = (3'd6);
  assign y8 = (3'd1);
  assign y9 = (2'd1);
  assign y10 = (({a2,a1}>(b2^p14))?((a2<b1)!=$signed({b4})):((&(a3^~b2))<(~|(~^b1))));
  assign y11 = ($unsigned({2{({a1,b5}|{a0,b3,b4})}}));
  assign y12 = (~&{3{((!b2)||{4{a2}})}});
  assign y13 = (^((^{(^{(~|p13)}),(+{2{p5}})})^~({{1{b0}},(~p7),(~|p12)}>>(~|{{b4,p14}}))));
  assign y14 = (((p13|p8)+(5'd2 * p8))?{{3{p15}},{3{p5}}}:(5'd2 * (-p14)));
  assign y15 = ((a4+a3)>$signed((~&a5)));
  assign y16 = {$unsigned(a5),(4'd2 * a0)};
  assign y17 = (|p2);
endmodule
