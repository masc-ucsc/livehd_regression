module expression_00246(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((4'sd4)^~(5'd16))+{4{(-4'sd4)}}),{3{{2{(-2'sd1)}}}},{1{((~|(5'd27))<=((3'd5)>>>(5'sd2)))}}};
  localparam [4:0] p1 = (+(({4{(-5'sd14)}}||((2'd3)?(5'd8):(3'd0)))?(((5'd28)|(-5'sd6))+((2'sd0)>>>(2'sd0))):(((4'sd3)?(3'd0):(2'd3))<<<((5'd11)>>(-2'sd1)))));
  localparam [5:0] p2 = {(!{2{((5'sd9)!=(3'sd3))}})};
  localparam signed [3:0] p3 = {3{{(!(-2'sd0))}}};
  localparam signed [4:0] p4 = ((2'd3)<<(4'sd2));
  localparam signed [5:0] p5 = {(((3'd2)>(5'd28))===(^(4'd14))),((5'd0)?(5'd22):(2'd2))};
  localparam [3:0] p6 = (~((((-5'sd6)+(4'd0))^~{(-5'sd12)})!==((~|(5'sd7))!==((4'd10)<<(2'd1)))));
  localparam [4:0] p7 = (-4'sd1);
  localparam [5:0] p8 = ({((4'd12)>=(5'sd4)),((5'sd4)>>(5'd24))}<=({(-3'sd3),(5'sd7),(4'sd6)}&{{(-2'sd1),(5'd17)}}));
  localparam signed [3:0] p9 = {4{(4'd12)}};
  localparam signed [4:0] p10 = ((((2'd2)<<<(5'd31))?{(5'd21),(-3'sd1)}:((-5'sd1)?(5'd10):(-5'sd3)))?(2'd1):(((4'sd1)-(-5'sd2))?((5'd7)?(2'sd0):(5'd25)):((-3'sd2)?(-2'sd0):(5'd18))));
  localparam signed [5:0] p11 = ((~^({(2'd3)}^(3'd1)))|{{(5'd7)},(&(4'd4)),((5'd28)||(4'd12))});
  localparam [3:0] p12 = {4{(5'sd15)}};
  localparam [4:0] p13 = (((3'd2)+(2'd1))?((4'd5)>>>(-2'sd1)):(|((4'sd4)!==(2'd3))));
  localparam [5:0] p14 = (2'sd1);
  localparam signed [3:0] p15 = {{{(3'sd3)}}};
  localparam signed [4:0] p16 = ({1{(6'd2 * (2'd2))}}<((2'sd0)?(4'sd3):(-4'sd0)));
  localparam signed [5:0] p17 = (5'sd6);

  assign y0 = (^{(p14>>>p5),(|p3)});
  assign y1 = (p16?a3:b5);
  assign y2 = ($signed(((|(b3^~a5))^~((b5<p3)<(|p10))))>=((|{3{b1}})<(&(&{4{a0}}))));
  assign y3 = (|(~&((b0*p6)%p13)));
  assign y4 = (((^(b4?p3:p4)))?((p11)?(p9?a4:p0):$unsigned(b2)):(~|((^$unsigned((a4?b2:a2))))));
  assign y5 = (~&{3{(-{1{p4}})}});
  assign y6 = (&$signed(($unsigned(((^p16)%p3))?((p2>>>p11)?(p0?p6:p17):(^p2)):$signed((p5?p14:p5)))));
  assign y7 = {($unsigned(b3)?{a4,p10}:{p17,p2}),{(p12?a1:b5),(5'd19)},{{p13,p0,p7},(3'd7),(5'sd13)}};
  assign y8 = ((p2|p11)%a2);
  assign y9 = ((4'd11)==(6'd2 * (a1>=a2)));
  assign y10 = (5'sd14);
  assign y11 = (~&{(~(((a5===a1)?(a3^~b0):(+p5))<<<((p16<<p16)&&(4'd2 * p7))))});
  assign y12 = {{4{p9}},{(-2'sd1)}};
  assign y13 = (~&{2{((+p5)>{2{p2}})}});
  assign y14 = (+(2'd0));
  assign y15 = {2{({3{p13}}?(b2>=b2):({1{b1}}))}};
  assign y16 = ((~&(b2?p11:b4))^~(^(|(b5>>b0))));
  assign y17 = (+(((a3>>>b3)^~(a2==b5))^((b5!=b4)^~(p12-a1))));
endmodule
