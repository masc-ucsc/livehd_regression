module expression_00728(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{{4{{(5'sd11),(4'd1)}}}}};
  localparam [4:0] p1 = (-2'sd0);
  localparam [5:0] p2 = ({(-(2'd3))}?((5'd8)|(5'd1)):((2'd2)?(-2'sd0):(5'sd12)));
  localparam signed [3:0] p3 = ({(-5'sd12),((4'd5)?(-4'sd6):(4'sd7)),(5'd30)}<((4'd6)-((2'd0)&&(4'sd3))));
  localparam signed [4:0] p4 = {2{{4{((-2'sd0)<=(-3'sd0))}}}};
  localparam signed [5:0] p5 = {(((5'sd8)^~(5'd15))?{(-5'sd14),(4'd8),(4'd0)}:((-3'sd0)&&(-4'sd7)))};
  localparam [3:0] p6 = (!(5'sd3));
  localparam [4:0] p7 = ((-5'sd9)^(-3'sd3));
  localparam [5:0] p8 = (2'd2);
  localparam signed [3:0] p9 = (~^((2'd3)+(2'd2)));
  localparam signed [4:0] p10 = (((-2'sd0)&&(4'sd2))!=((-3'sd1)>(4'd2)));
  localparam signed [5:0] p11 = (((4'sd3)?(-3'sd2):(3'd3))?((2'd0)?(4'sd6):(3'd4)):{1{((2'd2)>>>(-3'sd0))}});
  localparam [3:0] p12 = {{(~&(4'd14)),(!(2'sd1))}};
  localparam [4:0] p13 = {((4'd14)>>>(4'd0))};
  localparam [5:0] p14 = ((((2'd2)?(3'd2):(5'sd11))?(~&(4'd6)):((2'd1)?(3'd3):(-4'sd0)))&(|((5'd21)?(5'd10):(5'd29))));
  localparam signed [3:0] p15 = ((~^(3'd0))|(!(2'd0)));
  localparam signed [4:0] p16 = ({(-(3'sd3)),{(2'd3),(-2'sd0),(4'sd7)},(!(4'sd1))}==(^(((-3'sd1)!=(5'd30))|((4'd10)?(5'sd11):(3'sd0)))));
  localparam signed [5:0] p17 = (((2'd2)==(2'd1))||((4'd11)+(2'd2)));

  assign y0 = (&(p10&&b4));
  assign y1 = (p9?p14:p11);
  assign y2 = (5'sd8);
  assign y3 = {b3};
  assign y4 = (((a2?b1:b0)?(a3?a4:b1):(5'd22))!==((b3!==b4)!=(4'd1)));
  assign y5 = ({2{{3{b0}}}}>>>{4{(a2==a4)}});
  assign y6 = (5'd2 * (5'd13));
  assign y7 = {2{b0}};
  assign y8 = (&{(!({{b4},{a5,a4,a0}}===(|(4'd0))))});
  assign y9 = ((a0|a3)>>(~^(|a5)));
  assign y10 = {(-(5'd29))};
  assign y11 = (((p7>>>p15)?(|p8):(p17?p15:p17))>>>((p15&&p8)^~(&(p11^~p2))));
  assign y12 = {{$signed((p3?p17:b5)),($signed(p2)),{p13,p8,b3}}};
  assign y13 = ({3{{1{(b5==b2)}}}}>>>({1{({1{p4}}<={4{a1}})}}||({4{p10}}^~{2{a4}})));
  assign y14 = {3{((-p15)<<(-a5))}};
  assign y15 = {1{(|(!{2{((&(&b2))?(2'd3):{2{b0}})}}))}};
  assign y16 = (-5'sd11);
  assign y17 = (~(-p7));
endmodule
