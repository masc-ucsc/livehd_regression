module expression_00695(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(4'd8));
  localparam [4:0] p1 = (-{((-(3'd5))<=((2'd2)?(-4'sd4):(3'sd3)))});
  localparam [5:0] p2 = ((((3'd7)+(-5'sd5))<((3'd6)===(5'd22)))>={1{{3{(5'd2 * (2'd0))}}}});
  localparam signed [3:0] p3 = (&{1{(3'sd0)}});
  localparam signed [4:0] p4 = ((5'd5)!==(-2'sd0));
  localparam signed [5:0] p5 = (((2'd0)|(4'd15))?((-5'sd12)&&(2'd2)):((-4'sd1)<(2'sd0)));
  localparam [3:0] p6 = (-5'sd5);
  localparam [4:0] p7 = ((((4'd2)==(3'd4))^((5'd1)<<<(-4'sd1)))==((~{2{(3'sd2)}})|((2'd2)>>>(3'd1))));
  localparam [5:0] p8 = ({{2{(3'sd1)}},((5'd24)>>>(4'd1)),((3'd7)?(3'sd1):(4'd13))}-({2{{(5'd6),(2'd1),(-4'sd7)}}}<={((5'd30)<=(5'sd13)),{(-3'sd0)}}));
  localparam signed [3:0] p9 = (~^(|(~&(|(|(^(~&(5'd20))))))));
  localparam signed [4:0] p10 = (({((-5'sd1)&(2'sd1)),((5'd9)|(-3'sd2))}==={{(~|(5'sd15))}})||{((4'd0)>>(5'd12)),(^((4'd4)|(2'd0))),{((-4'sd3)&(2'd2))}});
  localparam signed [5:0] p11 = (((2'sd1)?(^(4'sd6)):(^(3'd3)))?(!((2'd0)?(5'd27):(2'd2))):(((-5'sd0)?(2'sd1):(5'd0))+((3'sd3)?(-2'sd1):(5'sd13))));
  localparam [3:0] p12 = (^(-4'sd3));
  localparam [4:0] p13 = ((3'd1)^~{((4'sd1)?(5'd31):(3'd1)),((5'd0)>>>(2'sd1))});
  localparam [5:0] p14 = (-((((-2'sd1)&&(2'd1))|(~^(~(-2'sd1))))^(~|(&(~&(&{(2'd3),(5'd26),(3'd4)}))))));
  localparam signed [3:0] p15 = (6'd2 * ((3'd7)&&(5'd30)));
  localparam signed [4:0] p16 = (^(5'd2 * ((4'd7)<=(4'd13))));
  localparam signed [5:0] p17 = (&(~|(|(((|(5'd6))!==(~|(-5'sd3)))?((4'd5)?(4'd15):(4'd9)):((2'd0)?(3'sd2):(4'sd3))))));

  assign y0 = ((((a0|p1)+{1{a3}})&&{3{b0}})<=(!({4{p4}}&&(a0-b0))));
  assign y1 = (a0?p8:p11);
  assign y2 = (2'd0);
  assign y3 = (-{2{(~&{2{(!(p13?p17:p2))}})}});
  assign y4 = (((b3?b0:p13)?(b1>>b1):(^(~^b5)))^~(|{(~b1),{b2},(-b4)}));
  assign y5 = {1{{{4{p3}},(~^$signed({p3,b4,b5}))}}};
  assign y6 = (p8?b2:a5);
  assign y7 = {$signed((~&(p6+a3))),{p12,a5,p6},$unsigned($signed({p1,a2}))};
  assign y8 = {(^(((4'd13)-{(2'sd0)})<<(~|(|(3'd1)))))};
  assign y9 = (p7>>>p15);
  assign y10 = (4'd6);
  assign y11 = ((~^(+(($unsigned(p13)?(p13/a3):(p7))?((p17?p12:b5)?(a4?b0:b1):(a1&b2)):((~|a3)?(p14/p4):(&b5))))));
  assign y12 = (^(2'd0));
  assign y13 = (b0?b5:a4);
  assign y14 = (5'd2 * (b1<<<p8));
  assign y15 = $signed(((p15>>p8)<(|b4)));
  assign y16 = (4'sd0);
  assign y17 = (|(({a4,a3}^(p13>>a3))<<{{p16,b3,b5},(+(b4|p10))}));
endmodule
