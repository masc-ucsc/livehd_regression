module expression_00157(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(~(~&{(2'd3),(-3'sd2)})));
  localparam [4:0] p1 = (5'd2 * (~(|(5'd0))));
  localparam [5:0] p2 = {1{{2{(5'd26)}}}};
  localparam signed [3:0] p3 = (6'd2 * {2{(2'd3)}});
  localparam signed [4:0] p4 = (~^{4{((-3'sd1)>>>(5'sd5))}});
  localparam signed [5:0] p5 = (4'sd5);
  localparam [3:0] p6 = (((-4'sd4)<(5'd19))?((-4'sd1)!=(5'd3)):((5'sd12)*(5'd26)));
  localparam [4:0] p7 = {3{(5'd2 * (4'd4))}};
  localparam [5:0] p8 = (~((&(2'd0))<(4'd5)));
  localparam signed [3:0] p9 = {(-3'sd3),(3'sd2)};
  localparam signed [4:0] p10 = (((-4'sd2)<<<(-4'sd3))?((-2'sd0)?(3'd6):(5'd5)):((4'd9)?(-3'sd0):(3'd4)));
  localparam signed [5:0] p11 = (~&(!(~&(~&(|(~|{{3{(2'sd0)}},{(5'd9),(2'd3),(-3'sd0)}}))))));
  localparam [3:0] p12 = (~&(+(!(|(-4'sd0)))));
  localparam [4:0] p13 = (~&(4'd14));
  localparam [5:0] p14 = {3{(-(~^(&(-3'sd3))))}};
  localparam signed [3:0] p15 = ((2'sd1)||(3'd6));
  localparam signed [4:0] p16 = {(((3'd1)>=(3'd6))<<<((-5'sd2)^~(-4'sd6))),{((2'sd1)<=(4'd8)),((2'sd0)-(2'sd1)),{(5'd28)}}};
  localparam signed [5:0] p17 = (|(3'd1));

  assign y0 = (((+((a2?b1:a1)&$unsigned(b1)))<((a4^a0)===(b2>=a1))));
  assign y1 = {1{((p4?p13:b2)?(a0<<<b2):{1{p4}})}};
  assign y2 = ($signed(((2'd1)<<(a4!=b1))));
  assign y3 = (~(~&{1{({1{(~^$unsigned({4{a2}}))}})}}));
  assign y4 = (-3'sd0);
  assign y5 = (~^{(~^{(|p15),(+p7),(&p6)}),(2'sd1),(|{(~|a4),(p7==b0),(|a0)})});
  assign y6 = (+b1);
  assign y7 = (((&((a3*a4)))<=(~|(p6==a0)))^((a4<<<b4)%a1));
  assign y8 = ((&{2{{4{p14}}}})<(^(-{3{(!(5'sd1))}})));
  assign y9 = (^($unsigned((b0>=b3))===(4'd0)));
  assign y10 = (~|($signed((4'd7))));
  assign y11 = ((-((b0===a3)!=={3{a0}}))<=($signed(a0)?(p1?a1:p5):{2{a4}}));
  assign y12 = $signed((|((~^(&(2'd2))))));
  assign y13 = $unsigned((~|{2{{2{p13}}}}));
  assign y14 = ((~&(~^p8))?(p13?p17:p11):{p9,p9,p9});
  assign y15 = $unsigned(((((b1?b3:a4)<$unsigned(b2))|((a4)||(b1+b3)))===(((b2)<(b2|b0))&&(a4?a4:a1))));
  assign y16 = ((((!b4))?(&(-b0)):(b5?p10:p2)));
  assign y17 = (4'd4);
endmodule
