module expression_00449(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((!{4{(2'd1)}})?{2{(5'd23)}}:((-3'sd2)?(5'sd15):(-2'sd1)));
  localparam [4:0] p1 = ((~|((3'd1)|(3'd6)))/(2'd3));
  localparam [5:0] p2 = ({1{(4'd13)}}^~((5'sd2)&(2'sd0)));
  localparam signed [3:0] p3 = ((~((5'd27)|(4'd4)))/(-5'sd13));
  localparam signed [4:0] p4 = ((((5'd22)<<(5'sd0))&&((-3'sd1)-(2'd2)))?(4'd2 * (5'd9)):(-3'sd1));
  localparam signed [5:0] p5 = (~&((4'd11)?(((2'd2)<<(-3'sd1))<<((5'd2)>>(5'sd15))):(~^{1{(~|(&(3'd7)))}})));
  localparam [3:0] p6 = ((((-2'sd0)?(3'd5):(2'd2))?((3'd0)?(-2'sd0):(5'd11)):((5'd18)?(-4'sd6):(5'd16)))?(((2'd1)?(5'd21):(4'd9))?((2'sd1)?(-3'sd0):(-5'sd3)):((5'd6)?(4'd15):(2'd0))):(((2'd2)?(-2'sd0):(2'd2))?((5'sd15)?(3'sd0):(2'd1)):((-4'sd0)?(3'sd3):(4'd8))));
  localparam [4:0] p7 = ((3'd7)?(4'sd5):(5'd26));
  localparam [5:0] p8 = ((((-4'sd3)==(-3'sd0))>{1{(3'sd0)}})>>>{3{((5'd4)<=(5'd7))}});
  localparam signed [3:0] p9 = ((-5'sd1)?(5'd6):(4'd9));
  localparam signed [4:0] p10 = ((((4'sd0)>(-3'sd0))<={1{(3'sd3)}})<(((4'sd7)^(-4'sd1))?(4'sd0):((-2'sd1)?(2'd0):(3'sd0))));
  localparam signed [5:0] p11 = (4'd2 * ((5'd14)?(4'd15):(2'd2)));
  localparam [3:0] p12 = ((((5'sd4)>>>(2'sd0))^((-3'sd2)/(2'd0)))>=(((3'd5)<(4'sd4))^~((2'd0)||(2'd2))));
  localparam [4:0] p13 = {{((-3'sd3)^~(3'd2)),(3'd6),{1{(5'd19)}}},({4{(3'd6)}}||(-4'sd6))};
  localparam [5:0] p14 = {(({3{(5'd5)}}&{3{(5'sd6)}})&(((4'd1)===(-5'sd5))-{(3'sd1),(-5'sd4),(2'd2)}))};
  localparam signed [3:0] p15 = {4{(-((-3'sd2)>>(2'd3)))}};
  localparam signed [4:0] p16 = {2{{2{{1{(3'sd2)}}}}}};
  localparam signed [5:0] p17 = (((4'sd7)<<(4'd12))!={(3'd2),(2'd1),(5'sd4)});

  assign y0 = (((^(a0*b1))<<(5'd25))-(2'd1));
  assign y1 = (((2'd2)||((a0^p16)^(a5*b2)))^(-5'sd5));
  assign y2 = {3{{3{(b4||b3)}}}};
  assign y3 = (((p6!=p14)>(p4<=p5))?(~&((p10^~p2)/p3)):(&(~(~(p1-p14)))));
  assign y4 = {(a5||a2),{p11,p0},(a0!==b1)};
  assign y5 = ({1{(((5'd2 * p2))^~{(b5===b2)})}}+({3{p5}}?(p7>p8):(p9<<<p10)));
  assign y6 = (({3{(b3||b0)}}<<<{4{(a0>b0)}}));
  assign y7 = {1{$unsigned($signed(p8))}};
  assign y8 = (!{1{{(((b4?a1:b1)?(^a0):{4{a1}})?{(p13?b3:p9),{a0,p15}}:{{b1,b1,b4},(|b4),(-a3)})}}});
  assign y9 = (((a3>>p5)|(3'd0))-(2'd2));
  assign y10 = ((+{2{((+p7)>>>(p0&b5))}})!=((|({4{a1}}!==(a1!=a0)))<<(^(4'd2 * (^p8)))));
  assign y11 = ((&((~&(&(b5^a0)))||(~|(b1==b0))))!=(((~^a0)&&(b5>>>b1))<<<((a5||p15)>=(~&p7))));
  assign y12 = (($unsigned({(4'd2)})-({(p3<=p5)}>>(p5<=p13))));
  assign y13 = ((b5!==a5)^(~|p16));
  assign y14 = (((((4'd5)+(^p10))||{1{($unsigned(p12)^~(p11<p17))}})));
  assign y15 = (^(|(5'd11)));
  assign y16 = (^({b0,p3,p9}?(+(p1?b4:p10)):{2{p11}}));
  assign y17 = (((!p6))|{(p11?b4:p4)});
endmodule
