module expression_00996(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd1);
  localparam [4:0] p1 = {(!(~(&(2'sd1)))),{(^(~(4'sd4)))},(~&(+{(-2'sd0),(3'sd2),(-5'sd0)}))};
  localparam [5:0] p2 = {1{{2{{2{((-4'sd2)<=(3'd7))}}}}}};
  localparam signed [3:0] p3 = (((4'sd6)>=(3'd4))<=(^(3'sd3)));
  localparam signed [4:0] p4 = (3'd1);
  localparam signed [5:0] p5 = ((&{{(-2'sd1),(-4'sd3),(2'sd0)}})?(&((4'sd2)?(-4'sd3):(-3'sd0))):(~&((5'sd9)?(5'd9):(2'sd0))));
  localparam [3:0] p6 = {((~{(4'sd1),(3'sd0),(-5'sd13)})>((2'sd1)==(-5'sd10))),(((3'd6)<(2'd0))>>(~^((-3'sd0)-(2'd0))))};
  localparam [4:0] p7 = (^(((3'sd3)&&(5'd22))<<(5'd24)));
  localparam [5:0] p8 = ((4'd10)?{4{(3'd5)}}:((4'd12)=={1{(2'd1)}}));
  localparam signed [3:0] p9 = (((4'd3)?(3'sd1):(4'd10))==={2{(2'd2)}});
  localparam signed [4:0] p10 = (&({3{(~(4'sd5))}}?{2{((-5'sd8)||(3'd4))}}:(((-4'sd4)?(5'sd1):(4'd15))+((2'd3)<<(4'sd5)))));
  localparam signed [5:0] p11 = (({(-3'sd1),(4'd5),(-2'sd1)}||{(4'sd7),(-2'sd0)})-{((2'sd0)^(4'd14)),((-3'sd2)-(-2'sd1))});
  localparam [3:0] p12 = {3{((2'd1)?(4'd9):(5'd13))}};
  localparam [4:0] p13 = (|(-4'sd1));
  localparam [5:0] p14 = ((((3'd5)|(4'd11))===((3'd5)<<(2'd0)))^~{3{((5'sd15)-(5'd19))}});
  localparam signed [3:0] p15 = (^({((-4'sd0)==(-3'sd3)),(~(&(-3'sd2)))}===({4{(2'd2)}}==={(-4'sd1),(3'd2)})));
  localparam signed [4:0] p16 = (6'd2 * ((3'd5)&(5'd27)));
  localparam signed [5:0] p17 = (5'sd0);

  assign y0 = (b5?p17:b0);
  assign y1 = ((3'd6)?{(b3|a3),(a4>>b5)}:(5'd14));
  assign y2 = {(b0^~a4)};
  assign y3 = (((!(b1===a5))/b1)<<<(((b3*a4)||(b3%b1))>>>((~|b4)+(a0%p14))));
  assign y4 = (~|(&(&(|((-({p4}<<(p2!=p8)))^(&(~&{b1,b4,p3})))))));
  assign y5 = {1{({{4{p6}}}?((b3?p5:p3)>>>(p14>>>p15)):{(5'd9),(4'sd4)})}};
  assign y6 = {({1{{(p3<p15)}}}?$signed((p2?b2:p4)):{(^p17),(p14>p0)})};
  assign y7 = (!$unsigned({{b3,b0},{b4,p17},(a3>>b5)}));
  assign y8 = ((p1%b4)|(p0^~b5));
  assign y9 = (&(((p15||p16)>=(b4&&p8))>>>(-(6'd2 * (+(p13==a0))))));
  assign y10 = (~|(~^((2'd0)==((-((a5===b3)%b5))))));
  assign y11 = {(3'd4)};
  assign y12 = $unsigned(((((~b5)*(~&p1))==(~|(b3^p4)))>$unsigned(($signed((~$unsigned(b5)))^((p4<<<a1))))));
  assign y13 = {(~&(5'sd0))};
  assign y14 = {(|(+({(^b2),{3{b4}}}!=={(^b5),(~|a5)})))};
  assign y15 = {3{{2{{p17,p11}}}}};
  assign y16 = (!({p5,p11,b2}?{p16,b2}:(!p17)));
  assign y17 = ((4'd2 * (b0^p0))-(&((!((a5%p15)<=(p11-p14))))));
endmodule
