module expression_00754(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{((-5'sd13)+(-2'sd1))}};
  localparam [4:0] p1 = ((5'd2)<=(5'sd14));
  localparam [5:0] p2 = (~&((|((2'd0)||(4'd14)))?((4'd9)!=(2'sd1)):(+(|(-5'sd11)))));
  localparam signed [3:0] p3 = (({(-3'sd0),(-5'sd7),(5'sd14)}^((4'd0)>>>(3'd0)))===(~&(4'd2 * {((2'd0)|(4'd14))})));
  localparam signed [4:0] p4 = (-(|((3'd2)%(-5'sd12))));
  localparam signed [5:0] p5 = (((-2'sd0)^~(-5'sd14))<<<((5'd18)<<(-4'sd5)));
  localparam [3:0] p6 = (((+(2'd2))&&{(-3'sd2),(2'd1),(4'd9)})?({(4'd6)}^((5'd19)>>(3'sd2))):(|((4'sd4)?(4'd2):(5'sd3))));
  localparam [4:0] p7 = (|(~^(2'd1)));
  localparam [5:0] p8 = ((^(-(2'd3)))<(-4'sd5));
  localparam signed [3:0] p9 = (~^(&(3'd6)));
  localparam signed [4:0] p10 = ({1{((-3'sd2)?(-2'sd1):(-2'sd0))}}?((2'sd0)?(-3'sd1):(2'sd1)):(5'd15));
  localparam signed [5:0] p11 = {(3'sd3),((4'd3)^(2'sd1))};
  localparam [3:0] p12 = {((((5'sd13)!=(4'sd1))<=((2'sd0)|(-2'sd0)))>=(~|((4'd7)?(3'd7):(5'sd6))))};
  localparam [4:0] p13 = (~&(4'sd4));
  localparam [5:0] p14 = (-5'sd5);
  localparam signed [3:0] p15 = (((3'd7)?(3'd2):(5'd11))!=(((-4'sd3)>>(3'sd1))==((-5'sd11)-(2'sd1))));
  localparam signed [4:0] p16 = ((5'sd5)?(5'sd9):(-2'sd0));
  localparam signed [5:0] p17 = {4{{4{(2'd3)}}}};

  assign y0 = {((-a1)>>(5'sd3)),(^(!(p3>>p6))),{1{(&(!(~p1)))}}};
  assign y1 = (+((~^{$signed((p3)),(~|(p0<p8))})<((6'd2 * p0)>>(!(+p3)))));
  assign y2 = ((5'sd8)!==({a3,b3}-(-4'sd6)));
  assign y3 = (5'd2 * (^(-b1)));
  assign y4 = ((a1|b0)/p14);
  assign y5 = (((b5<b5)<<{a1,a5})||((a5>a5)|(b5-b2)));
  assign y6 = (~(2'sd0));
  assign y7 = ((p8>b4)<(-2'sd0));
  assign y8 = ($signed(((p9?a1:p10)<<$unsigned(p5)))?((p11?b1:p0)?(b3<<p11):(p14)):$unsigned($unsigned(((b1&p2)<(p7?a2:a1)))));
  assign y9 = {{(4'd13),(4'd9),(b3!=a5)}};
  assign y10 = (($signed((&$unsigned(p16)))>{2{(p17>>>p10)}})>(((p10^~a3)<<{{p3}})));
  assign y11 = (p0>>p5);
  assign y12 = ({{1{{(b0||b3),{a5,b2},$signed($unsigned(p8))}}},((~{3{p17}})?(a5?b5:p1):(a2?a3:b5))});
  assign y13 = {p4,p1};
  assign y14 = {(p10<=p13),{a0,b0,b3},$unsigned((~&b3))};
  assign y15 = ((&(p13?p10:p10))?((a0===a0)>>>{4{b0}}):{1{(~^{1{{4{p9}}}})}});
  assign y16 = (~(({(a1),{b2,b5,b5}}<<<{a0,a1,a4})!={($signed((a3?b4:a5))?(a3>=b5):(b5?b3:b5))}));
  assign y17 = {3{($unsigned((~b2))<<<{4{a5}})}};
endmodule
