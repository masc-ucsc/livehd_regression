module expression_00279(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd0);
  localparam [4:0] p1 = (|((3'sd1)?(-2'sd0):(5'sd0)));
  localparam [5:0] p2 = {((3'd4)==(5'd16)),(3'd2),(!(3'd5))};
  localparam signed [3:0] p3 = {1{(((2'sd1)===((2'sd1)&(3'd5)))>=({4{(3'd7)}}>=((4'sd3)<(4'sd0))))}};
  localparam signed [4:0] p4 = (+(&(~&{2{({4{(4'd0)}}&&((3'd4)>=(-5'sd2)))}})));
  localparam signed [5:0] p5 = {1{(5'sd12)}};
  localparam [3:0] p6 = (2'd0);
  localparam [4:0] p7 = (-(5'sd11));
  localparam [5:0] p8 = ((((-5'sd8)?(2'sd1):(-3'sd0))<={2{(-2'sd1)}})>=((2'd3)?((3'd6)?(2'd3):(4'sd6)):(~|(4'sd3))));
  localparam signed [3:0] p9 = {4{(2'sd0)}};
  localparam signed [4:0] p10 = (!((-4'sd4)<<<(5'd4)));
  localparam signed [5:0] p11 = {3{(~&(((5'd29)<<(2'd0))^~{(3'sd2),(5'sd1)}))}};
  localparam [3:0] p12 = {4{(2'd2)}};
  localparam [4:0] p13 = {3{(4'd1)}};
  localparam [5:0] p14 = (((3'd4)>>(2'd3))?{(4'sd0),(-4'sd0),(-2'sd0)}:(-4'sd0));
  localparam signed [3:0] p15 = (((3'd6)?(5'd12):(5'd13))?((4'd5)>(3'd1)):((2'sd0)?(-4'sd3):(3'd1)));
  localparam signed [4:0] p16 = (((2'd0)^~(3'd4))?((-4'sd4)&&(3'sd3)):((2'd1)&(2'd2)));
  localparam signed [5:0] p17 = (-((5'sd12)?(4'd0):(4'sd1)));

  assign y0 = (5'sd10);
  assign y1 = (~&p10);
  assign y2 = ((4'd8)+((~^$unsigned((3'sd2)))===((^b1)^(b2>>a4))));
  assign y3 = $unsigned({1{$signed((({1{$unsigned({3{b3}})}}!==({3{b1}}-$unsigned(a5)))>>>($signed((p4<<p12))<={2{{3{a1}}}})))}});
  assign y4 = (+(&(^(4'd1))));
  assign y5 = {2{p6}};
  assign y6 = ((((a2>b0)<={1{b4}})>>>$signed(((p11)>(a5))))>>(4'd2 * $unsigned($unsigned(b3))));
  assign y7 = {2{{3{b0}}}};
  assign y8 = (-((~{(~^p12)})?{(^p16),(&p3)}:((p5?b3:b0)||(p3<<b4))));
  assign y9 = (a0>>p17);
  assign y10 = {{(~|p5),(p8+p12),(p11<<b1)},(-((|b1)===(b1||b1))),(~^{4{p5}})};
  assign y11 = (~|(|((~^p15)!=(^p13))));
  assign y12 = $signed(($signed(((~(p8&p17))<=(p14?p5:p4)))));
  assign y13 = {{(b1<<<a5),{a3,b3,p4}},(2'sd1)};
  assign y14 = (((a3?b0:p10)<{{3{b1}},(&b3)}));
  assign y15 = (-(~&((p6&&b2)^(p1|p2))));
  assign y16 = (+(~^{(b4==b3),(a5&b5),(!(3'd6))}));
  assign y17 = ((((b5&&p4)+{p13,b0,p4})!=((p9>>p0)!=(p2||a1)))-{{{{{(p15-p12),{p10,p11,p15},(p3|p9)}}}}});
endmodule
