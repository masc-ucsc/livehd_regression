module expression_00621(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-2'sd0)<=(((2'd1)!=(3'sd1))&((2'sd0)==(4'sd2))));
  localparam [4:0] p1 = (4'sd6);
  localparam [5:0] p2 = (+(-4'sd2));
  localparam signed [3:0] p3 = (6'd2 * {{(3'd3)}});
  localparam signed [4:0] p4 = ((|((5'd19)?(3'd6):(3'd4)))|((-2'sd1)?(3'd6):(4'sd2)));
  localparam signed [5:0] p5 = (|(&(+(+{4{((5'sd9)?(-3'sd1):(2'd1))}}))));
  localparam [3:0] p6 = (~^{(~|((5'sd5)?(-5'sd11):(-4'sd6))),{(3'd0),(4'd8)}});
  localparam [4:0] p7 = (^{4{(5'd11)}});
  localparam [5:0] p8 = ((-4'sd6)<(3'd3));
  localparam signed [3:0] p9 = (~&(+(~&(-4'sd0))));
  localparam signed [4:0] p10 = ((((-5'sd8)==(4'd13))?((-4'sd6)<<(-4'sd4)):{(3'd6),(2'd2),(3'd1)})+({(-5'sd2)}?(3'd4):(4'd14)));
  localparam signed [5:0] p11 = (4'd15);
  localparam [3:0] p12 = {(~|(-{(-5'sd7),{(-4'sd2),(2'd0),(4'd4)}}))};
  localparam [4:0] p13 = ((4'sd2)/(-4'sd7));
  localparam [5:0] p14 = (!(((5'd30)?(4'sd1):(5'd8))?((4'sd1)?(3'd6):(4'd10)):{3{(5'sd5)}}));
  localparam signed [3:0] p15 = (^{((4'd10)?(2'd3):(-4'sd3)),((4'd15)?(5'd25):(4'sd3)),{(-5'sd5),(4'd9)}});
  localparam signed [4:0] p16 = (-4'sd2);
  localparam signed [5:0] p17 = {4{((2'd1)?(3'sd3):(2'd2))}};

  assign y0 = {1{{((p11)>>>(~b0)),{1{({p6,p11}=={4{p1}})}}}}};
  assign y1 = {2{(b1!==b3)}};
  assign y2 = (3'd3);
  assign y3 = $signed((~&(!{4{((-p13)^(p4^~p3))}})));
  assign y4 = (3'd6);
  assign y5 = (b0|b5);
  assign y6 = ($signed((~^(p10?p3:p4)))?(p16?p8:p6):$signed({4{p7}}));
  assign y7 = ($signed({2{(a4|a1)}})&($signed(a0)!==(b3>a1)));
  assign y8 = {{1{($signed(((p6^b0)>>>(b3==b3))))}},(^(^({a4,b4,a1}>>(~^(6'd2 * b0)))))};
  assign y9 = {(~^{{b1},(~|p10),$unsigned(a5)})};
  assign y10 = {2{((b2?b2:p8)?(p13?p17:a0):(a5))}};
  assign y11 = (&(~^{(~|(5'sd0)),(~|{p7,a5}),(b1?p3:a2)}));
  assign y12 = (((&(p8?p14:b0))-(p11?p7:p16))&(~(~&((p0&&p12)!=(p7<<p1)))));
  assign y13 = ((((a1-a5)>>(a4+b2))+((b3*a0)!==(~&a4)))>>>(~|(+(5'd2 * (b2||p1)))));
  assign y14 = (({b5,a0}!==(-b0))^(&(5'd10)));
  assign y15 = {((b3===b5)+(b4<=b5)),(4'd2 * {(b1^a0)}),(!(+(+{p17,p5})))};
  assign y16 = $signed((2'sd1));
  assign y17 = ((!(b1<<p0))^{{(^b1)}});
endmodule
