module expression_00512(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{3{((4'd4)>>>(2'd2))}});
  localparam [4:0] p1 = {3{(2'd2)}};
  localparam [5:0] p2 = (~|(~&(-5'sd3)));
  localparam signed [3:0] p3 = {(3'd0)};
  localparam signed [4:0] p4 = ((|{1{{1{(^(!{3{(3'd1)}}))}}}})&&(((5'sd4)&&(4'sd1))<=((5'd7)>=(4'd6))));
  localparam signed [5:0] p5 = (3'd6);
  localparam [3:0] p6 = ((~|((3'd3)?(2'sd1):(3'd3)))?((4'sd3)?(5'd26):(5'd8)):(5'sd4));
  localparam [4:0] p7 = ((((-4'sd3)?(5'd21):(2'd1))>(+(4'd14)))!=(((2'd0)?(-2'sd1):(2'd1))-((2'd0)||(-4'sd1))));
  localparam [5:0] p8 = {4{{4{(3'd2)}}}};
  localparam signed [3:0] p9 = (+((!{3{(5'd8)}})?(^(^((-5'sd15)?(4'sd2):(-5'sd13)))):(^{4{(2'd1)}})));
  localparam signed [4:0] p10 = (|(~^(((~((-5'sd1)*(4'd5)))&(~^((-3'sd2)-(5'd17))))!==((~(!(5'd6)))==(!((4'd3)^(4'd14)))))));
  localparam signed [5:0] p11 = ((((4'sd2)===(3'd3))^((4'd1)||(-3'sd2)))+(((2'd1)||(2'd3))%(-4'sd0)));
  localparam [3:0] p12 = (+((2'sd0)?((-2'sd0)|(-5'sd10)):((5'd0)>>(2'd3))));
  localparam [4:0] p13 = (((3'sd2)||(2'd1))===((3'sd2)===(-4'sd4)));
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = ({1{((-3'sd2)!=(3'd3))}}?{1{((3'd0)<<<(3'sd1))}}:(((-5'sd12)?(3'd6):(3'd1))<<<((2'sd1)?(5'd12):(-4'sd2))));
  localparam signed [4:0] p16 = (((((2'sd0)<<<(4'sd4))&((2'd3)>=(-2'sd1)))|((!(3'd1))||((2'd0)!==(4'd3))))<=((((-3'sd0)^~(5'sd15))<<(6'd2 * (2'd2)))>>(+((5'd12)^(3'sd0)))));
  localparam signed [5:0] p17 = ({(((4'sd6)?(2'd2):(4'sd3))?((-2'sd1)?(-2'sd1):(-3'sd3)):((-4'sd5)?(3'sd0):(4'sd1)))}&&(((4'sd6)||(4'sd0))?((-3'sd0)?(4'sd6):(4'd9)):((5'd31)!=(4'd14))));

  assign y0 = {{{{({a5,b5,b3}?(p3?a5:b1):{b2,p15}),{{b4,p17,p9},{b1},(a3?b0:a5)},{{b5,b5,a0},(b5?b1:p15)}}}}};
  assign y1 = (b2&&b0);
  assign y2 = ({4{(+(p8<b5))}});
  assign y3 = (a5===a0);
  assign y4 = ({1{{4{a0}}}});
  assign y5 = {1{{1{({1{{1{((5'd12)==={3{a1}})}}}}<<(-3'sd3))}}}};
  assign y6 = ({4{b4}}<=({p14,a0}&&(+a4)));
  assign y7 = (((~&(a5===a4))<<(a3==a1))^($signed(($signed((b3>=b3))))));
  assign y8 = (|(+(~($signed({4{p6}})>>>({{2{b4}}}==(&{p14,a1}))))));
  assign y9 = {2{p4}};
  assign y10 = (3'd3);
  assign y11 = ((-4'sd1));
  assign y12 = (2'd2);
  assign y13 = {({b0,a0}&&{a1,b4}),{1{{2{a1}}}}};
  assign y14 = (^(~^(-(~&($unsigned({$unsigned((p0+a1)),{(~|p12)}})&(!(~&(-4'sd7))))))));
  assign y15 = ((-((p16)!=$unsigned(p10))));
  assign y16 = ({p17,b4}==(p16||a4));
  assign y17 = ((p4?p17:p0)?(~p13):(a1+a2));
endmodule
