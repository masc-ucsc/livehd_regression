module expression_00366(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(&(-5'sd13))}};
  localparam [4:0] p1 = {(-4'sd1),(-4'sd7),(-2'sd0)};
  localparam [5:0] p2 = {2{((!(4'd3))=={4{(2'd0)}})}};
  localparam signed [3:0] p3 = {4{(3'd2)}};
  localparam signed [4:0] p4 = (3'd1);
  localparam signed [5:0] p5 = (({(4'd12),(3'd7)}?((4'sd5)>>(4'd4)):((2'sd1)?(5'sd4):(-4'sd1)))&&(((-4'sd5)!=(2'sd0))^~((-4'sd4)!==(-3'sd2))));
  localparam [3:0] p6 = (~^(&(+(!(!(|(~(&(!(3'd0))))))))));
  localparam [4:0] p7 = ((((2'd0)-(-4'sd7))<={(4'd7),(5'd12),(3'sd0)})===(((4'd8)<=(4'd11))>>>((-2'sd1)?(4'd7):(4'sd3))));
  localparam [5:0] p8 = (~^{{3{{(2'd3)}}},({(2'sd0)}?{(5'd12)}:{(2'd2)})});
  localparam signed [3:0] p9 = ((-4'sd3)<=(2'sd1));
  localparam signed [4:0] p10 = (-(((~&(2'sd0))>(4'd2 * (2'd0)))?((|(4'd3))?((3'd4)?(3'd4):(5'sd6)):((4'd0)<<(3'sd0))):(((3'd1)^~(5'sd9))?((2'sd1)<<(3'd4)):(~(3'sd1)))));
  localparam signed [5:0] p11 = ((~^(3'd2))?((3'd1)&(2'd1)):((3'd5)-(4'sd0)));
  localparam [3:0] p12 = ((3'sd2)>>(3'd2));
  localparam [4:0] p13 = (4'd12);
  localparam [5:0] p14 = (-4'sd2);
  localparam signed [3:0] p15 = (~&(-((5'd28)?(3'd4):(5'sd3))));
  localparam signed [4:0] p16 = {(^(3'd1))};
  localparam signed [5:0] p17 = (-((4'd3)?(5'd21):(5'd13)));

  assign y0 = {1{{1{{1{{1{a4}}}}}}}};
  assign y1 = (3'd7);
  assign y2 = $unsigned((2'sd0));
  assign y3 = (|{((|({a3,a4,p14}<=(b3&&p14)))?{{b3,a4},{b0},{a2,b5,a1}}:(~&{(b2&b5),{a5,b3}}))});
  assign y4 = ({4{p1}}?(2'd2):(4'sd3));
  assign y5 = (4'd0);
  assign y6 = {4{(a3)}};
  assign y7 = ((p5||p17)*(!(a4!=p3)));
  assign y8 = (+(~(((&b0)&(-p16))<=((a0==p1)<<(b4>a0)))));
  assign y9 = (!(!{(-4'sd2)}));
  assign y10 = (((b4==p7)%p7)+(((b2/a3)<=(b4&b3))>>>((b1*b2)<(b0>>b5))));
  assign y11 = ({2{p14}}<=(4'd0));
  assign y12 = (a5?b1:a4);
  assign y13 = {{2{(((p15?p15:b2)-(5'd18))>>{4{a2}})}}};
  assign y14 = (((b1<b1)<(b0||a4))>((a2+b0)==(a2||a3)));
  assign y15 = (~&(((p13>b0)||(p7+p3))&(&(5'sd6))));
  assign y16 = (6'd2 * (p12?b1:p13));
  assign y17 = (((-b3)<=(3'd2))!==((&b0)!=(b1>b5)));
endmodule
