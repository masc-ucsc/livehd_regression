module expression_00258(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~({1{{1{(3'd1)}}}}<{2{(2'sd1)}}));
  localparam [4:0] p1 = {1{((((5'sd5)?(5'd20):(3'd5))?{4{(-4'sd4)}}:{(5'd19)})!=(((4'd15)-(5'd15))>((5'd18)&(2'd0))))}};
  localparam [5:0] p2 = (^(|(+((|(~|(-2'sd0)))>=((3'd0)<<(4'sd3))))));
  localparam signed [3:0] p3 = (|(&(3'd6)));
  localparam signed [4:0] p4 = (5'd27);
  localparam signed [5:0] p5 = (5'sd5);
  localparam [3:0] p6 = (~|(-(^(|(~(&(+(+(&(~^(3'sd1)))))))))));
  localparam [4:0] p7 = {1{((4'd1)-((3'd5)?(2'd2):(-5'sd6)))}};
  localparam [5:0] p8 = {{(5'd31),(5'd2),(3'sd0)},((2'd3)===(5'd2))};
  localparam signed [3:0] p9 = (|((~(|{((~(4'sd4))>={(2'd2),(4'd6),(2'd1)})}))<<(&(!((~&(3'sd0))&&(3'd5))))));
  localparam signed [4:0] p10 = (&(-(((5'd19)?(5'd14):(-3'sd2))?((^(4'd10))<<(~(5'd19))):{2{(~^(3'sd1))}})));
  localparam signed [5:0] p11 = {4{{1{(5'sd15)}}}};
  localparam [3:0] p12 = (((4'sd3)==(-2'sd1))?(|(-2'sd0)):((3'sd0)?(-2'sd0):(3'sd0)));
  localparam [4:0] p13 = (((5'd13)^(-2'sd1))?((3'sd1)?(5'sd0):(5'd27)):{(3'sd2),(2'sd1),(2'd1)});
  localparam [5:0] p14 = (&((5'd4)!=(^(5'd7))));
  localparam signed [3:0] p15 = (~^(~&(^(-(4'd1)))));
  localparam signed [4:0] p16 = (-2'sd1);
  localparam signed [5:0] p17 = {(2'sd1)};

  assign y0 = (~((~|((~|((~&p3)))<(~$signed((p9<<<p4)))))));
  assign y1 = {3{(^a4)}};
  assign y2 = {({(a1!==a0),{3{p13}}}<<{(^{p8})}),{3{{3{p12}}}}};
  assign y3 = {{(5'd10),(a2?p5:p2)},(2'd0)};
  assign y4 = {2{(~(!($signed(p0)==(p16!=p0))))}};
  assign y5 = (2'd0);
  assign y6 = ((p0?p2:p10)?(3'd0):{2{p9}});
  assign y7 = (~$unsigned((((b2||a2)===(b2>b1))>>>(|(~^{p1,b5})))));
  assign y8 = (!{2{{4{(^a3)}}}});
  assign y9 = {{b0,p9,a5},(a1?a5:a5)};
  assign y10 = (-(-2'sd0));
  assign y11 = (|(2'd3));
  assign y12 = (-(p16?b2:p9));
  assign y13 = (+{a4,p16,p8});
  assign y14 = ({(~|(p8>>>p2)),(p1<<p15),(p1<<<p6)}<<{({p14}>={p0,p2,p15}),{(^{p12,p13,p14})}});
  assign y15 = {((-(~p10))!=(5'd2 * p2)),({p3,p10,p14}=={(~p2)})};
  assign y16 = (4'd2 * (2'd3));
  assign y17 = (4'd14);
endmodule
