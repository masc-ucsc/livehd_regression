module expression_00802(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd3)?(-2'sd1):((-2'sd0)&(2'sd1)));
  localparam [4:0] p1 = (+({{((4'd9)<(-5'sd0))}}===(-((-5'sd4)<<(3'd1)))));
  localparam [5:0] p2 = ((((5'd18)?(4'sd2):(5'sd8))?((2'd2)===(2'sd0)):(+(3'd2)))&&{{(-3'sd1),(4'd8)},(~(4'd3)),((3'd7)?(5'd12):(4'd2))});
  localparam signed [3:0] p3 = ((4'd8)?(3'd7):((3'd4)||(5'd20)));
  localparam signed [4:0] p4 = (4'd5);
  localparam signed [5:0] p5 = (((3'sd2)^~(4'd12))&&((3'd5)>=(3'd3)));
  localparam [3:0] p6 = ((((-3'sd3)?(3'd2):(3'd0))?((4'd8)?(5'd1):(5'd6)):((2'd2)?(2'd3):(-2'sd1)))?{3{((2'd1)<<<(3'd4))}}:(4'sd1));
  localparam [4:0] p7 = (((-4'sd1)>>>(5'd31))<((3'd3)>>(3'sd3)));
  localparam [5:0] p8 = {3{(~&{2{(2'd3)}})}};
  localparam signed [3:0] p9 = ((((4'd7)?(5'd2):(2'sd1))>>((4'd11)<<<(4'sd4)))|{4{(-(3'd5))}});
  localparam signed [4:0] p10 = {2{{2{{1{((3'd5)<<<(3'd4))}}}}}};
  localparam signed [5:0] p11 = (!(~(!(4'd8))));
  localparam [3:0] p12 = (!{(-(~&(~&(|((4'd0)?(2'd3):(-2'sd0)))))),(~&(~{4{(3'd4)}}))});
  localparam [4:0] p13 = {3{(2'd3)}};
  localparam [5:0] p14 = ((-(-((~&((3'd5)>>(3'd6)))>={((5'd22)-(-3'sd3))})))+(~&(-{{(2'd3),(3'sd0)},(~(&(5'sd0)))})));
  localparam signed [3:0] p15 = {1{(4'd2 * {2{(3'd3)}})}};
  localparam signed [4:0] p16 = (~&((4'sd6)||(3'd6)));
  localparam signed [5:0] p17 = (|(-(~^(~(-(~|(&(!(|(~^(~&(4'd13))))))))))));

  assign y0 = (+((a3?a4:p13)?{1{(4'd4)}}:{3{p6}}));
  assign y1 = $unsigned(($signed({2{(p2|p9)}})<{(p0<<<p14),(~^p10),(p8^~p17)}));
  assign y2 = ((|(((a3|p6)<=(~|p10))|{(~|b5),(a5&&a0)}))|($signed((a0+a4))===(^{(~|a0)})));
  assign y3 = (~&((a2!==a5)?(-b4):(|p9)));
  assign y4 = $unsigned(((p16/p10)));
  assign y5 = {2{((-a0)?{p16,p0}:{p13})}};
  assign y6 = (3'd7);
  assign y7 = (4'd3);
  assign y8 = (|((a4-a4)<=(!(a2))));
  assign y9 = ((p6?b2:p14)*(~(p2>>>p17)));
  assign y10 = (((5'd12)<=(+a5))===((a0<b0)==(b4!=b1)));
  assign y11 = ((+(-5'sd10)));
  assign y12 = (({3{$unsigned(p0)}}-{1{(p11?p14:p13)}})==(((p8?p11:b1)?(p6?p4:b4):(p8!=p14))==((p12?b1:p16)?(p11?p14:p11):(p3==p17))));
  assign y13 = ($unsigned(b5)<=(a0^p5));
  assign y14 = ((b0?p5:a1)?(b3?a1:a5):(~|b4));
  assign y15 = {(~^{2{{(2'd1),(2'sd0)}}}),{{1{{(a5?b4:p9),(+(p1?p15:p15))}}}}};
  assign y16 = $signed($signed($unsigned($unsigned((~|(|(~(^$unsigned(((~|$signed((~^p6)))))))))))));
  assign y17 = ((b0-a5)<<<(a2<a3));
endmodule
