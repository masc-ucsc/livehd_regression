module expression_00685(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd3)>>(5'd5));
  localparam [4:0] p1 = (~(((~^(3'd0))+((4'd2)-(3'sd2)))^(!(((-3'sd1)!==(3'd1))>=(&(-4'sd3))))));
  localparam [5:0] p2 = (({(5'd29),(3'sd2),(3'd6)}>>((2'sd0)!==(2'd3)))<{3{{2{(5'sd13)}}}});
  localparam signed [3:0] p3 = (^{4{(~&(2'sd1))}});
  localparam signed [4:0] p4 = ((((2'sd1)>(-3'sd2))>>>((-2'sd0)^(2'd2)))^((+((-3'sd0)&&(5'd2)))+((4'd9)&&(4'sd7))));
  localparam signed [5:0] p5 = (~&{(-4'sd5),(5'sd6),(3'sd1)});
  localparam [3:0] p6 = (~|(~&(!(~|((2'sd1)!==(-3'sd3))))));
  localparam [4:0] p7 = (({(4'd14)}<((3'd1)===(2'd1)))==(((4'd0)<<(3'sd1))=={(4'sd7),(4'd14),(3'sd3)}));
  localparam [5:0] p8 = {(2'd1),(5'd5),(-3'sd0)};
  localparam signed [3:0] p9 = (((2'd3)==(2'd3))>={(3'd0),(5'd0),(3'd0)});
  localparam signed [4:0] p10 = {(((-4'sd6)?(5'd6):(3'd1))?{(-4'sd7),(4'd5),(3'd3)}:{(-5'sd5),(3'd5)}),(((-4'sd6)?(4'sd5):(-5'sd0))?((4'd10)?(4'sd2):(4'd13)):((4'd4)?(-4'sd2):(-5'sd1)))};
  localparam signed [5:0] p11 = (~|(((-(!(5'd7)))>>>((5'sd15)^~(2'd3)))!=(~((~^(~^(3'sd1)))-(-((2'sd1)===(5'd10)))))));
  localparam [3:0] p12 = (~&{{(~({2{(-5'sd4)}}&&{(4'sd5),(4'd6)}))}});
  localparam [4:0] p13 = (-2'sd0);
  localparam [5:0] p14 = ((4'sd6)&&(3'd5));
  localparam signed [3:0] p15 = ((|((~|(-5'sd3))/(4'd4)))?((4'd2 * (3'd1))/(2'sd1)):((^(4'd4))?((3'sd0)==(2'd0)):((-3'sd1)&(3'sd0))));
  localparam signed [4:0] p16 = ((((4'd10)?(2'd3):(3'd6))<={{(4'd13)}})>>>(((-2'sd0)?(5'd19):(3'd5))?(~(2'd0)):(~&(5'd10))));
  localparam signed [5:0] p17 = ((((-2'sd0)>>(5'd3))===((2'd3)<<<(3'sd1)))<<(((-5'sd11)>>>(-3'sd3))^((-5'sd3)!==(5'sd1))));

  assign y0 = (4'd8);
  assign y1 = (|(!(b1>>p13)));
  assign y2 = (-(((b0||a5)^(5'd25))<<<((b0&a1)>(a0===a1))));
  assign y3 = (b2&&b5);
  assign y4 = {$signed((({((+(~a5))>(b0!=a2))}))),((+((p10!=p17)>=$signed(a3)))^~(~^(+(a1&&b4))))};
  assign y5 = $unsigned((((p9?a0:a4)<=$unsigned(b0))?{1{(p1?p2:p6)}}:{((a2?b4:a0))}));
  assign y6 = ((&(b3>=b4))>(a2>>b0));
  assign y7 = (|(~|(b2?p0:p3)));
  assign y8 = (({(p6==a0),(a0?p14:p12),(p8?p11:p6)}<{$signed(a4),{1{a2}},(p5>>p12)}));
  assign y9 = (p15<p11);
  assign y10 = {((b5^p7)<<<(~|p3)),{(a5?p15:a4),(b3-a1)},$signed(((p10+a4)))};
  assign y11 = (&(~|(~^(-({3{(&(p9<=a0))}}&((~|(~|(~b3)))^(~|(~^(a3===a4)))))))));
  assign y12 = (3'sd3);
  assign y13 = ((+(&(b5<b4)))!==((b5||b0)-(-2'sd0)));
  assign y14 = (~|(p3>>>a5));
  assign y15 = ($signed((p12-b3))*((p10>=p2)));
  assign y16 = (3'd2);
  assign y17 = {(~^(a2===b0)),((b4>>>a3)===(!b4)),((+a1)<<{a4,a1})};
endmodule
