module expression_00374(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd4)?(~&((3'sd3)?(5'd31):(2'sd1))):(((3'd3)||(-4'sd1))?(5'd1):(^(2'd1))));
  localparam [4:0] p1 = (((3'sd1)>>(4'd2))/(2'd1));
  localparam [5:0] p2 = ((((3'd4)?(4'd12):(4'sd2))!=={((-5'sd13)<(3'sd1))})<(-2'sd1));
  localparam signed [3:0] p3 = ({3{(~(2'd3))}}<<<{((2'd0)?(3'd3):(4'd8)),(-(5'sd15))});
  localparam signed [4:0] p4 = (|{{({{(3'sd0)}}^~{(^(3'd3))}),(((-3'sd3)>(-2'sd0))&(&((4'd15)!==(2'd3))))}});
  localparam signed [5:0] p5 = {2{{3{((2'd2)!==(2'd3))}}}};
  localparam [3:0] p6 = (~^(((~^(5'd28))<((-3'sd3)?(4'd10):(2'd3)))>>>(((3'd4)!==(4'sd7))^((-4'sd5)&&(3'sd2)))));
  localparam [4:0] p7 = {1{{2{(~|({4{(-3'sd0)}}>>((4'sd0)?(2'd2):(5'd12))))}}}};
  localparam [5:0] p8 = (~^(((3'd3)-(3'd1))?(|((-2'sd0)^(5'd20))):((5'd12)||(2'sd1))));
  localparam signed [3:0] p9 = {{(4'sd4),(&{2{(5'd29)}}),(~&(4'd5))}};
  localparam signed [4:0] p10 = (-2'sd0);
  localparam signed [5:0] p11 = {3{{(2'd0),(3'sd2)}}};
  localparam [3:0] p12 = (((5'sd5)&(5'd6))?((5'sd1)===(-4'sd3)):((4'sd4)?(4'sd7):(2'sd1)));
  localparam [4:0] p13 = ((3'sd3)?(-4'sd7):(3'd1));
  localparam [5:0] p14 = (4'd2 * ((5'd5)<<<(4'd0)));
  localparam signed [3:0] p15 = (&((4'sd1)/(4'd13)));
  localparam signed [4:0] p16 = (~&{1{((~|(((3'sd0)?(-3'sd0):(-4'sd7))|(!(4'd8))))|(-((-3'sd3)?(-2'sd1):(4'd11))))}});
  localparam signed [5:0] p17 = (~|{4{((3'sd2)<(-2'sd0))}});

  assign y0 = $unsigned($signed($signed(($signed($signed((4'd5)))))));
  assign y1 = ((a0+p16)%b0);
  assign y2 = (~|(&(-($signed(((&p8)))?((b3>=b0)!=={b0,b4}):((a2===b4)&&(~^p3))))));
  assign y3 = $signed({4{$signed(p11)}});
  assign y4 = (4'd4);
  assign y5 = ((!(|p15))<<<(p5?p4:p15));
  assign y6 = ($unsigned((a0!==b4))?(({1{p14}})):{4{a2}});
  assign y7 = $signed({3{(({3{p8}}>>>$unsigned(p17)))}});
  assign y8 = (~(+(~&(-{{((b4?p2:a4)?(p13?a0:p6):{2{(p0?p14:p4)}})}}))));
  assign y9 = (^$unsigned(({(5'd2 * (-(p13-p12)))}>=(((~&(+p6))+{p13,p7,p17})))));
  assign y10 = (3'd3);
  assign y11 = (!(b3-p14));
  assign y12 = ((^{b1,b2,a2})===(!(b2!=b4)));
  assign y13 = (4'd5);
  assign y14 = {4{((4'd11)<(p16==p12))}};
  assign y15 = (~{4{{4{p16}}}});
  assign y16 = ((~(~|(!((~^p7)<(b1===a1)))))>=((!(b1|b3))!==(~(5'd2 * a1))));
  assign y17 = (p5^~p9);
endmodule
