module expression_00906(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((&(+(2'sd1)))<<<((2'd2)?(2'd2):(4'd15)))<=((-5'sd3)<<((4'sd0)?(3'd3):(4'd14))));
  localparam [4:0] p1 = (({2{(2'sd1)}}-((2'sd0)==(-3'sd3)))>>(+((6'd2 * (4'd7))?{2{(5'd1)}}:{3{(-5'sd9)}})));
  localparam [5:0] p2 = (3'sd0);
  localparam signed [3:0] p3 = {(-4'sd3)};
  localparam signed [4:0] p4 = (3'sd1);
  localparam signed [5:0] p5 = (|((((3'sd3)^(3'sd3))===((5'd10)?(-4'sd2):(4'sd3)))&(-(5'sd13))));
  localparam [3:0] p6 = ((3'd5)||(-3'sd3));
  localparam [4:0] p7 = (4'd3);
  localparam [5:0] p8 = ((^(~^{3{(~&(3'sd1))}}))>(^(5'd2 * (&(~|(3'd0))))));
  localparam signed [3:0] p9 = (&(5'sd7));
  localparam signed [4:0] p10 = (2'd2);
  localparam signed [5:0] p11 = {4{{(5'd22),(-3'sd1),(2'd1)}}};
  localparam [3:0] p12 = ((~(-(3'd2)))?(~&((-3'sd0)?(-3'sd0):(2'sd1))):(~|(-(2'd0))));
  localparam [4:0] p13 = ((~((~^(4'sd3))>>((3'd7)?(2'd2):(5'sd5))))?(((3'd4)>>>(5'd16))?(&(2'd0)):((2'd1)?(3'sd0):(-4'sd4))):(~(|((4'd8)&&(3'd7)))));
  localparam [5:0] p14 = (&(^(|(!(5'sd0)))));
  localparam signed [3:0] p15 = (((5'd11)>>(2'd3))<<<{2{(5'd10)}});
  localparam signed [4:0] p16 = ((5'd18)?(5'd25):(-5'sd9));
  localparam signed [5:0] p17 = {((4'sd3)?(2'd1):(-4'sd6))};

  assign y0 = ((p3?p2:b1)>>(p13?p4:b2));
  assign y1 = {{(~{1{(b3-a2)}}),(-2'sd0)},(~^(^(5'd31)))};
  assign y2 = (((~&{(~&(|a5)),(^$unsigned(a0)),(~&(p15<<b4))})||{$unsigned((~^{(!$unsigned(p10)),$signed($unsigned(a3))}))}));
  assign y3 = {2{b4}};
  assign y4 = (p15<=a1);
  assign y5 = ((p2>>>p2)<(&p13));
  assign y6 = (~(~|$signed((a0===a2))));
  assign y7 = (((&(~&p6))>>((-p12)))<={1{$unsigned((-(&(~&a0))))}});
  assign y8 = (-3'sd3);
  assign y9 = (a2-b0);
  assign y10 = (^(-2'sd0));
  assign y11 = {3{(5'sd5)}};
  assign y12 = (~^(-(~|(5'd12))));
  assign y13 = (4'd4);
  assign y14 = ((p9<<p14)&{b2,p5});
  assign y15 = (!((p14|p8)>>(b1*p0)));
  assign y16 = (((p16>b4)>=(b1||p17))?((b0<<b5)!=(b4<b2)):((p6?a0:a4)^~(a0>>b2)));
  assign y17 = (p7&&a5);
endmodule
