module expression_00229(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd2 * ((4'd8)&(2'd2)));
  localparam [4:0] p1 = (~^((~(+({3{(4'sd6)}}&((5'd9)&(5'd15)))))||(~(~&({2{(2'd0)}}<((4'sd5)||(2'd0)))))));
  localparam [5:0] p2 = (4'sd6);
  localparam signed [3:0] p3 = (~^({(5'd29),(4'd1),(4'sd0)}|(^{(3'd4),(2'd1)})));
  localparam signed [4:0] p4 = (~(~&(((4'd2)<(5'sd11))<((4'd12)===(2'd2)))));
  localparam signed [5:0] p5 = (-(~|(!(6'd2 * (~^((5'd29)+(4'd9)))))));
  localparam [3:0] p6 = ((5'd3)!==(-2'sd1));
  localparam [4:0] p7 = (^(&((((3'd6)|(-5'sd15))+((2'd3)!=(5'sd3)))&&((~^(2'sd0))^(!(2'd3))))));
  localparam [5:0] p8 = (-4'sd6);
  localparam signed [3:0] p9 = {2{{2{((-3'sd2)>(4'd7))}}}};
  localparam signed [4:0] p10 = (^(~^(2'd2)));
  localparam signed [5:0] p11 = (~|(((5'd10)===(-4'sd0))^~(|(2'd0))));
  localparam [3:0] p12 = ({1{(-2'sd1)}}?(~&(4'd1)):((5'd19)?(3'd2):(2'd2)));
  localparam [4:0] p13 = {((^{({(-4'sd3),(4'd1)}>>(^(5'd10)))})>>((|(^(-5'sd3)))+{2{(3'd6)}}))};
  localparam [5:0] p14 = {{(-2'sd1),(5'sd6)},(~&(5'sd7))};
  localparam signed [3:0] p15 = ((5'd7)>>(2'sd0));
  localparam signed [4:0] p16 = (-(5'd28));
  localparam signed [5:0] p17 = ((((5'd31)%(-5'sd8))?((4'sd0)!==(-4'sd5)):((5'sd4)^~(3'd2)))!=(((5'd17)&(2'sd1))===((4'd6)?(4'sd5):(4'd3))));

  assign y0 = (3'd1);
  assign y1 = (p1|a0);
  assign y2 = (((-(-2'sd1))>=((4'd2 * a2)-(~p16)))==((|(~^(6'd2 * p8)))>=(-3'sd2)));
  assign y3 = {2{{3{p4}}}};
  assign y4 = (p3?p13:p0);
  assign y5 = (((a3&b4)!==(b2&b2))>>{2{(-p15)}});
  assign y6 = ((b4===a5)%b5);
  assign y7 = (5'd15);
  assign y8 = {2{(-(~|{3{(p1>p3)}}))}};
  assign y9 = ({(~p2),(b2?b0:a2),(~^a5)}?{(-3'sd1),(2'd1)}:{(2'd0),(p8?a5:a3),(~^p14)});
  assign y10 = ((((a3?a5:b2)+(a1&a2))!==(b1?b5:b2))^~(((6'd2 * p7)<<<(p3^~p17))||((5'd2 * p12)-(p3||b1))));
  assign y11 = (a2>>>a3);
  assign y12 = (4'd15);
  assign y13 = (((~(-3'sd1))>>{3{(+a0)}})<({(p14&p4),(-4'sd6)}<<<((p5>>p13)-(~|p4))));
  assign y14 = (((($signed((~|b5))?(~(^a2)):(b3-a4))>>>(+((a5>>>b0)?(b5&a2):(p6?b1:a0))))));
  assign y15 = (-(~|({{(~b5),{p8},(|a5)}}^{(p6>=p15),(~^p1),{p16}})));
  assign y16 = {{3{(~&(~{{3{a0}}}))}}};
  assign y17 = (((b1<=b4)>=(b5^~b4))-((b4<p5)|(p15>>>b2)));
endmodule
