module expression_00800(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~|(-3'sd1))<((3'd5)||(2'd2)));
  localparam [4:0] p1 = (~^{1{(~|(~|{(-4'sd5),(3'd1)}))}});
  localparam [5:0] p2 = (((4'sd3)-(2'sd0))?(~&(3'd5)):((4'sd1)?(-5'sd13):(2'sd1)));
  localparam signed [3:0] p3 = (({1{(2'd0)}}^((3'd3)>>(2'sd0)))?((3'd7)?(2'sd1):(2'sd1)):({(-2'sd1)}===(+(5'd29))));
  localparam signed [4:0] p4 = (5'd12);
  localparam signed [5:0] p5 = {{(-4'sd4),(-5'sd13),(4'd4)}};
  localparam [3:0] p6 = ({{(-3'sd0),(3'd3),(2'sd0)}}?(~^{(~|{(-5'sd4),(-2'sd1),(-2'sd0)})}):(^((4'd5)?(5'sd3):(-2'sd0))));
  localparam [4:0] p7 = ((~&(((-3'sd2)+(-2'sd1))>=(~&((2'sd1)^(4'd4)))))<=(~&(^((^(!(-3'sd0)))-(~^((3'd1)|(2'sd1)))))));
  localparam [5:0] p8 = {4{({1{(2'd1)}}<<<((-4'sd1)>(5'sd10)))}};
  localparam signed [3:0] p9 = (~&(+(+(+(^(~&((~|{4{(5'd10)}})?((3'd0)?(5'd13):(-3'sd3)):((3'd1)?(-5'sd6):(2'd1)))))))));
  localparam signed [4:0] p10 = ((2'd3)^~(2'sd1));
  localparam signed [5:0] p11 = {2{(|(-(!(2'd1))))}};
  localparam [3:0] p12 = (4'd7);
  localparam [4:0] p13 = ((((5'd9)>>(2'd2))<((-3'sd3)||(3'd4)))<<<((-(-4'sd3))^~(!(2'd1))));
  localparam [5:0] p14 = (5'sd13);
  localparam signed [3:0] p15 = {2{((~&(5'd4))<=(~|(3'd4)))}};
  localparam signed [4:0] p16 = (3'd1);
  localparam signed [5:0] p17 = ((3'd2)>=(5'd31));

  assign y0 = (^(5'sd13));
  assign y1 = (((p13?p8:a2)>>>$signed(p0))>=((p9)>>(~p2)));
  assign y2 = (6'd2 * {p6,a1});
  assign y3 = (^(~(((b4?a3:a1)?(b2?a3:a5):(~^(a4!==b0)))>=((5'd2 * {3{a0}})===((b4!==a0)&&(a3<=a1))))));
  assign y4 = {2{(-{2{{3{p2}}}})}};
  assign y5 = ($unsigned({2{(5'd8)}})===(5'sd3));
  assign y6 = {(~p1),(p5?p9:p0)};
  assign y7 = {{{{{p15,a4,b0}}},{{p16,b5},{p1}}},(({p4,b2}+(p15<=p8))<<({p1}?(p14?a2:p14):{a1,b4}))};
  assign y8 = (|(~&{3{{4{b0}}}}));
  assign y9 = (a5^~p0);
  assign y10 = ($unsigned({4{b0}})!=(a5<a3));
  assign y11 = (5'd20);
  assign y12 = $signed((~|(&$signed({({p8,p2,b4}<<<(~^(a4)))}))));
  assign y13 = ((((a5^~b3)!==(a5!=a1))>({3{p1}}>{p6}))!={(({p10,p12,p3}<=(p16|p8))<=((b1!==b4)>>>(-p3)))});
  assign y14 = ($unsigned((^a5))<(p5==b0));
  assign y15 = ((b5===b5)<=(p17&p11));
  assign y16 = {$unsigned({{a0,a2},$signed(b4),(a4)}),{{{a3},{a3,p5},$signed(p8)}},{$unsigned($unsigned(p11)),$signed($unsigned(b5))}};
  assign y17 = (&(~|p1));
endmodule
