module expression_00021(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd8);
  localparam [4:0] p1 = (+{1{(!(&{4{(3'd0)}}))}});
  localparam [5:0] p2 = (5'd11);
  localparam signed [3:0] p3 = (~|(~^(+(-{4{(~|(3'd5))}}))));
  localparam signed [4:0] p4 = (~^(((~(4'sd7))^~((3'd5)?(4'd10):(-3'sd0)))-((-(4'sd4))/(3'd3))));
  localparam signed [5:0] p5 = (~^{(~^({((2'd1)?(4'sd1):(2'sd1))}?((-2'sd0)?(5'd13):(5'sd3)):((4'd10)?(-2'sd0):(5'sd10))))});
  localparam [3:0] p6 = ((&(((-3'sd1)&(2'd0))!==(^((5'd12)>>>(5'd16)))))<<(((-2'sd0)&&(-5'sd8))<=(+((-3'sd3)<<(3'd3)))));
  localparam [4:0] p7 = (|{1{(|(+(6'd2 * (^(~^(5'd20))))))}});
  localparam [5:0] p8 = (((2'd0)?(-2'sd0):(-4'sd7))|(&((-3'sd0)?(3'd3):(4'sd3))));
  localparam signed [3:0] p9 = (~|(|(2'sd1)));
  localparam signed [4:0] p10 = ((3'd0)-(5'd19));
  localparam signed [5:0] p11 = {1{{(-4'sd0),(2'sd1),(2'd3)}}};
  localparam [3:0] p12 = ((((5'sd7)?(-5'sd9):(5'sd10))>>>((-5'sd1)<<(2'd0)))<<<(!{2{((2'd3)?(4'd12):(-5'sd1))}}));
  localparam [4:0] p13 = (!((3'd2)?(5'd28):(3'd4)));
  localparam [5:0] p14 = (~^(|(((2'd3)?(3'sd2):(2'd0))&&(~^((-2'sd0)==(-2'sd1))))));
  localparam signed [3:0] p15 = ((((5'sd6)?(3'sd1):(-5'sd2))<=(6'd2 * (5'd8)))||((!(3'sd3))>=(-(-2'sd0))));
  localparam signed [4:0] p16 = (((-2'sd1)?{3{(2'd0)}}:((-5'sd5)?(3'd7):(5'sd1)))!=({1{((-4'sd0)^(-5'sd4))}}===(-3'sd2)));
  localparam signed [5:0] p17 = (((-2'sd0)?(5'd20):(2'd1))?((4'd0)?(-5'sd4):(2'sd1)):((2'sd0)?(-3'sd2):(4'd13)));

  assign y0 = (2'sd0);
  assign y1 = ({2{$unsigned(p6)}});
  assign y2 = (3'd4);
  assign y3 = (p7==p5);
  assign y4 = ((a4?b4:a2)==(a4?b5:p8));
  assign y5 = ({{2{p9}},(p0!=p16),(2'd2)}^$unsigned(({3{p6}}^~{p14})));
  assign y6 = (5'd16);
  assign y7 = ({(p11|p7),(p9?p10:p17)}?({3{p10}}?{p14,p10}:{a1,p9}):{{3{b5}},(p10&&p1),(p6||p9)});
  assign y8 = ($signed((3'd1))===(4'd14));
  assign y9 = (~^(-(^(&(((~&(b2&&b2)))<<<(^{(4'sd4)}))))));
  assign y10 = (~^((~(-3'sd3))==((-(p11?b4:b2))%b5)));
  assign y11 = (!{(+(-{(~|(~&(|(~|(-p17)))))})),{{p5,p3,p4},(+{{p7,p2}})}});
  assign y12 = (~(5'sd8));
  assign y13 = (&(~|p14));
  assign y14 = (($unsigned($signed({p10,p10}))==(-((b1<b5)||(p12==a4)))));
  assign y15 = ((5'd17)^~((b2!==a0)+(p1%b5)));
  assign y16 = ($unsigned(p17)?(b3?b4:b0):(&p10));
  assign y17 = ({3{{2{$signed({2{p1}})}}}});
endmodule
