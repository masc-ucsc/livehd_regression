module expression_00731(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{({1{(~(((5'd10)?(-3'sd1):(3'sd3))<=((2'sd1)&(-4'sd3))))}}&({1{(|(-2'sd0))}}==((-3'sd2)+(3'sd2))))}};
  localparam [4:0] p1 = ((((4'd1)?(3'd2):(4'd10))>((2'd3)||(3'd0)))?(^((-5'sd10)?(-5'sd2):(-5'sd10))):(~((4'd7)-(3'd3))));
  localparam [5:0] p2 = ({{3{(3'd3)}},{(-3'sd2)}}&&{{1{{(4'd0),(2'd1)}}}});
  localparam signed [3:0] p3 = (|({((-3'sd0)?(-5'sd4):(-3'sd1)),(^(5'd4)),(~|(3'd1))}?(((3'd4)?(3'sd1):(4'sd3))?((2'd1)?(4'd8):(4'sd0)):{(5'd2),(3'd2),(3'd6)}):{2{((3'd0)?(-5'sd6):(-3'sd2))}}));
  localparam signed [4:0] p4 = ((~&(((5'd26)==(-3'sd1))?(5'd2 * (3'd6)):((4'd14)?(5'sd11):(-3'sd3))))-(((-2'sd0)?(4'd11):(-4'sd0))<={(5'sd7),(3'd5),(5'd6)}));
  localparam signed [5:0] p5 = {{(2'd2),(2'sd0)}};
  localparam [3:0] p6 = (((2'sd0)?(2'sd1):(3'd4))!=={(2'sd1),(4'd1),(2'sd1)});
  localparam [4:0] p7 = {3{((5'd14)<(2'sd0))}};
  localparam [5:0] p8 = {(~&{(3'sd0)})};
  localparam signed [3:0] p9 = ((((-2'sd0)<(3'd0))==((4'd6)<<<(3'd1)))<<<(((3'd2)>>(4'd14))==((5'd12)-(5'sd12))));
  localparam signed [4:0] p10 = (((4'd2)|(-2'sd0))<((3'd2)^~(3'd2)));
  localparam signed [5:0] p11 = (~(~^{2{(^(5'd30))}}));
  localparam [3:0] p12 = (+((~^(-2'sd1))=={3{(-3'sd3)}}));
  localparam [4:0] p13 = {(-3'sd3),(5'd5),(3'sd1)};
  localparam [5:0] p14 = ((-2'sd1)||((2'd2)-(4'd0)));
  localparam signed [3:0] p15 = {3{(2'd1)}};
  localparam signed [4:0] p16 = ((2'sd0)&&(-4'sd2));
  localparam signed [5:0] p17 = (((2'd2)==(5'd5))*(4'd12));

  assign y0 = {b5,a1,b4};
  assign y1 = (p17&&p0);
  assign y2 = $unsigned((+(&$signed((2'd3)))));
  assign y3 = ({(!(|({p15,a3,b3}))),{(|((b0<a1)<<<(~^a4)))},((b1^~p6)==(~&(p15==p13)))});
  assign y4 = (6'd2 * p13);
  assign y5 = $signed($unsigned({3{$signed(a3)}}));
  assign y6 = $signed((5'sd1));
  assign y7 = ({p14,p7}<<<(p4!=p15));
  assign y8 = (($signed((&(-2'sd0)))<{(a4),(3'd6)}));
  assign y9 = (~(!(&((&(4'd2 * (^b1)))==(&((~|p5)>=(p2|p4)))))));
  assign y10 = (p5?p16:p9);
  assign y11 = {2{p17}};
  assign y12 = (~|(-({3{(b4+a4)}}?$signed(((4'sd7)&&(p13>>>p10))):(-3'sd3))));
  assign y13 = ((((a4||a3)>=(~^a4))===((a2&&a0)|(b5<=a2)))<(~&(((b0&&b2)>>(b4>a2))!==(+(b5&&a5)))));
  assign y14 = (({4{p4}}-(~&a4))>=(((p7?p12:p16)^(p15?p3:a5))));
  assign y15 = (((a3&&p15)?(-5'sd2):(!p14))&(~((2'd2)?(p6^~b1):(-p9))));
  assign y16 = (~^p0);
  assign y17 = {3{{3{b5}}}};
endmodule
