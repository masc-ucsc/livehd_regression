module expression_00018(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{4{(5'd22)}}}};
  localparam [4:0] p1 = {4{((4'd1)==(2'sd1))}};
  localparam [5:0] p2 = {{(4'sd4),(4'sd3)},((4'd2)-(-4'sd4)),((-3'sd1)||(-3'sd2))};
  localparam signed [3:0] p3 = (((((5'd18)<<<(4'sd1))||(|(2'sd0)))<<<(~^(^((2'd0)&&(4'd2)))))<((^{1{((4'd12)===(-4'sd7))}})^~(-((-2'sd0)|(-2'sd1)))));
  localparam signed [4:0] p4 = ((((4'd9)&&(-4'sd0))^((5'd24)%(-4'sd4)))>=((6'd2 * (4'd10))*(3'd2)));
  localparam signed [5:0] p5 = ((((3'd2)>(5'sd15))<<(4'd2 * (5'd27)))>(((3'sd0)%(3'd4))^~((-2'sd1)>>>(2'sd0))));
  localparam [3:0] p6 = (((4'd0)?(2'd0):(2'd3))?(~|(5'sd12)):(4'sd7));
  localparam [4:0] p7 = ((-3'sd2)?(-4'sd3):(5'd22));
  localparam [5:0] p8 = {3{(!(4'd10))}};
  localparam signed [3:0] p9 = ((((5'sd9)^(5'd12))*((-2'sd1)^(2'd0)))-(((4'd8)>(2'd0))<((3'd2)!==(3'd6))));
  localparam signed [4:0] p10 = (-3'sd1);
  localparam signed [5:0] p11 = (~&(+(~^(~&{(2'd0)}))));
  localparam [3:0] p12 = {({((2'd2)?(-5'sd8):(2'sd1)),{(2'sd0)},{(5'd31)}}?(((-2'sd1)?(5'd23):(3'd5))?((5'sd0)?(4'd15):(-2'sd1)):((5'd6)?(5'd22):(3'd1))):{{(5'd10)},((4'sd1)?(-3'sd0):(4'd3))})};
  localparam [4:0] p13 = (3'd6);
  localparam [5:0] p14 = (~&(~^(-2'sd1)));
  localparam signed [3:0] p15 = ((3'd2)===((2'sd1)||(3'sd0)));
  localparam signed [4:0] p16 = (-(6'd2 * (+{(2'd1),(5'd9)})));
  localparam signed [5:0] p17 = (((4'sd6)==(-5'sd7))>=((2'd1)>=(-4'sd6)));

  assign y0 = $signed((({2{p15}}>(p11!=p1))&&{4{{2{b1}}}}));
  assign y1 = ((~|(^(-2'sd1)))^((a1?b5:a3)?(b3?a4:b5):(+(^p1))));
  assign y2 = (((-{p16,a5,p17})+(b2||p16))-((p12-a1)<(a5||b4)));
  assign y3 = (^(&(-(~|(~^$signed($signed((-((p2?a1:p2)?(p12):(p11?p3:p6))))))))));
  assign y4 = ({4{{4{a4}}}}?(-((p1?b0:p0)?(-5'sd12):(4'd12))):((~p1)?{1{p11}}:(!b0)));
  assign y5 = ({1{(4'd2 * {1{(p7||p14)}})}}||((p4?p0:p2)?(p2-p15):(a1===b1)));
  assign y6 = (3'd7);
  assign y7 = (^((-2'sd1)?(4'd14):(b4?p11:p2)));
  assign y8 = (4'd12);
  assign y9 = (!((((p10)>=(+p11))>>({p14,b4,p16}))&{3{(a4!==a3)}}));
  assign y10 = (b4>p0);
  assign y11 = (|{3{(p4>p13)}});
  assign y12 = {2{(&p9)}};
  assign y13 = {({p13,b1,p9}>(b1^~b1)),{1{{b5,b0,p12}}},({p13}>={4{a0}})};
  assign y14 = (-(&{(p7<<<p10),(p6<p0)}));
  assign y15 = ($unsigned(((a1?a1:b2)-(b2>>>b3)))>>>(-(((b1?b2:a4)==(-5'sd10)))));
  assign y16 = (p0>>p6);
  assign y17 = ({1{(p9<=a3)}}>((p2==p16)>>(p17&&p0)));
endmodule
