module expression_00084(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(2'd1),(5'd18)},((4'd2)>>>(2'sd1))};
  localparam [4:0] p1 = (4'd2 * ((4'd4)<=(5'd10)));
  localparam [5:0] p2 = {2{(((3'sd2)&&(3'd1))?{2{(2'd2)}}:(4'd3))}};
  localparam signed [3:0] p3 = (~|((+(((4'sd4)==(2'd3))|(^((4'sd0)<(-2'sd1)))))^~(((2'd2)&(3'd6))%(4'd5))));
  localparam signed [4:0] p4 = {((4'd3)==({(5'd22),(4'd15),(3'sd2)}<<<{((4'd7)>=(-2'sd0))}))};
  localparam signed [5:0] p5 = (~&(-3'sd3));
  localparam [3:0] p6 = {2{(2'sd0)}};
  localparam [4:0] p7 = (((4'sd7)?(2'd2):(4'd1))&((2'd1)?(-2'sd0):(4'sd5)));
  localparam [5:0] p8 = ((((-3'sd1)%(4'sd7))&((4'd15)^(3'd6)))==(((2'd1)!=(-4'sd0))-((5'd23)?(5'd15):(5'sd12))));
  localparam signed [3:0] p9 = {3{({4{(4'sd4)}}>{(3'd3),(4'sd3)})}};
  localparam signed [4:0] p10 = (5'sd0);
  localparam signed [5:0] p11 = (3'sd1);
  localparam [3:0] p12 = {{(2'd2),(-4'sd4),(3'd1)}};
  localparam [4:0] p13 = {2{(-4'sd3)}};
  localparam [5:0] p14 = {3{(-2'sd0)}};
  localparam signed [3:0] p15 = (~^(|(3'd0)));
  localparam signed [4:0] p16 = (3'd3);
  localparam signed [5:0] p17 = ((2'd3)?(2'd2):(3'd1));

  assign y0 = ((5'd11)<<((p11<<<p8)>>>(p11>a0)));
  assign y1 = (~^$signed((a4+p11)));
  assign y2 = (({b5,p17,a3}=={1{p14}})<<(+((p1>p10)<=(p15<<p9))));
  assign y3 = ({3{$signed($unsigned($unsigned(b5)))}});
  assign y4 = (~&({{p13,p4,p3}}<{p9,p4,p8}));
  assign y5 = {1{({(4'd2 * (p2>=p0)),{3{p8}}}&{1{({p4}?{4{b3}}:(p7?b4:p10))}})}};
  assign y6 = ($signed(p5)?(p12>>a1):(p0||p5));
  assign y7 = (|((~&$signed((!b3)))));
  assign y8 = (({a0}||{b5,a1,a3})!==((b4&&b4)==(a0||b5)));
  assign y9 = (((p9?b4:b1)+(5'd29))?((a2-a5)>(3'd2)):((b0>>a3)!=(p2?b3:b1)));
  assign y10 = {2{((~|(5'd15))?(p16?a1:p2):(^(5'd19)))}};
  assign y11 = {(~^$unsigned(b2)),(-3'sd2),(&(3'd4))};
  assign y12 = $signed((3'd7));
  assign y13 = (|((|p17)||{4{b3}}));
  assign y14 = ((((a5>=a0)|(b1!==a5))-({3{b0}}==(p13<<<b1)))&&{1{(((p17^~p6)&(a3|a2))<((a5&p6)^~(a3&a4)))}});
  assign y15 = {(+(p5||p12)),(-(a2<<b0)),(&(p17?b3:a5))};
  assign y16 = (~^{2{{1{$unsigned({2{a4}})}}}});
  assign y17 = ((a5?b4:b0)?$signed((a3<=b5)):{4{a0}});
endmodule
