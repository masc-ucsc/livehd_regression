module expression_00268(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~^(5'd1))>>>((5'sd5)&&(4'sd5)))>>>(((5'sd4)^~(-2'sd0))>>((4'd7)!==(5'sd0))));
  localparam [4:0] p1 = {2{{3{{2{(5'd0)}}}}}};
  localparam [5:0] p2 = {3{(4'd2)}};
  localparam signed [3:0] p3 = (~|(-5'sd3));
  localparam signed [4:0] p4 = {(((5'd5)?(3'sd3):(5'd16))?((2'd2)!==(4'd5)):{{(-3'sd2)}})};
  localparam signed [5:0] p5 = ((((5'd2)?(-4'sd0):(2'd2))>((-3'sd2)?(-4'sd1):(3'd5)))!=(((4'd5)^(5'sd10))+(5'd28)));
  localparam [3:0] p6 = ((4'd11)|(2'd3));
  localparam [4:0] p7 = {3{((-2'sd1)?(5'sd12):(-5'sd2))}};
  localparam [5:0] p8 = ((~&(~|(2'd2)))%(5'sd6));
  localparam signed [3:0] p9 = ((!(^(-5'sd9)))>((-2'sd1)>>>(2'd2)));
  localparam signed [4:0] p10 = {(2'sd0)};
  localparam signed [5:0] p11 = (((5'd1)/(5'd8))?((-2'sd1)-(-4'sd2)):((3'd0)?(4'd13):(-4'sd2)));
  localparam [3:0] p12 = {((~^{(2'sd1),(-2'sd0)})?(~|{(3'sd0),(-4'sd4)}):{1{{4{(5'sd6)}}}})};
  localparam [4:0] p13 = ({(2'd1),(4'd1),(4'sd1)}^{(-4'sd6)});
  localparam [5:0] p14 = (!{1{({{(5'd17),(3'd0),(4'sd2)}}||{4{(2'sd0)}})}});
  localparam signed [3:0] p15 = (((4'sd5)==(-2'sd1))||((-3'sd2)-(2'd0)));
  localparam signed [4:0] p16 = ({((2'd1)!==(-2'sd0)),{(3'd5),(5'd26),(5'sd14)},{(-4'sd7)}}||(((5'd28)+(-4'sd7))!==((4'd6)?(4'd4):(3'd4))));
  localparam signed [5:0] p17 = (-5'sd10);

  assign y0 = (4'd2 * (!{a2,b0}));
  assign y1 = ((p7?a1:p8)<<<(~&(a1&p7)));
  assign y2 = ((!((|(2'd1))!=(|(b3>=p12))))&&(~(((-3'sd2)||$unsigned(a1))+((p5|a2)^~(a3^~p11)))));
  assign y3 = {$signed(((4'd1)))};
  assign y4 = (5'd2 * (p7+p8));
  assign y5 = (4'd2 * (b2&p14));
  assign y6 = (((~^p15)?(a2?p8:p12):(5'd2 * p2))+(-((p4&&p0)<(p14<<p10))));
  assign y7 = (((-2'sd1)<{b1,b3,b1})?({a0}^~(p9)):((a5<<<p1)?(p10+p6):(5'd2 * p0)));
  assign y8 = ((4'd2 * {b0,a1})?(3'd1):((-2'sd1)>(a4<a5)));
  assign y9 = (^$unsigned({(~^{a5,a0}),(3'd6),(3'sd3)}));
  assign y10 = (~|{(p17>>>p5),(p13&p5),{3{p13}}});
  assign y11 = (|({4{(b3==a3)}}));
  assign y12 = {{{1{({(a2<<<a3)}^~({1{a5}}&{3{a1}}))}},({1{(a4^~p6)}}&&((b4>b4)>={2{b1}}))}};
  assign y13 = ((a3?p4:p8)?(5'd22):{2{(5'd29)}});
  assign y14 = (~(~$signed(($signed((~|((~^p2)<<<$signed(a0))))^$signed((~|(|((!p12)<=(^p14)))))))));
  assign y15 = {1{(p9?p7:p13)}};
  assign y16 = (!(p11>>>p15));
  assign y17 = (+p13);
endmodule
