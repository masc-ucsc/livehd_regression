module expression_00202(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd13);
  localparam [4:0] p1 = (~(3'd3));
  localparam [5:0] p2 = (((5'd4)?(-2'sd0):(4'd15))/(-4'sd6));
  localparam signed [3:0] p3 = {3{{2{(2'd3)}}}};
  localparam signed [4:0] p4 = (2'sd0);
  localparam signed [5:0] p5 = ((((5'sd12)>>>(3'd6))<{2{(-4'sd7)}})>{3{(4'd6)}});
  localparam [3:0] p6 = {{((-(5'd14))?((-3'sd3)?(3'd4):(3'd4)):((5'd17)>>(4'sd1))),(((3'sd1)?(5'd2):(5'sd0))^(~^(-5'sd11))),(((4'd12)-(2'd2))?((2'd0)!=(5'sd14)):((4'sd7)?(3'd4):(3'd1)))}};
  localparam [4:0] p7 = ((2'sd0)?(5'd7):(5'd3));
  localparam [5:0] p8 = {(~|(~&(2'd2)))};
  localparam signed [3:0] p9 = (3'd2);
  localparam signed [4:0] p10 = (~&(3'd0));
  localparam signed [5:0] p11 = ((-5'sd15)&&((!(3'sd3))?(3'sd1):((-2'sd0)?(5'd4):(4'sd0))));
  localparam [3:0] p12 = (^(~|((~|(|(2'sd1)))?((3'sd3)?(4'd9):(4'sd2)):((4'd7)?(3'sd3):(-5'sd4)))));
  localparam [4:0] p13 = ((((4'd12)|(5'd11))?((4'd6)!=(5'd13)):(-2'sd1))!=(((4'd5)>>(3'sd3))>((3'd6)&(-5'sd5))));
  localparam [5:0] p14 = (+({2{(4'sd7)}}?(~&(4'sd6)):{4{(2'd2)}}));
  localparam signed [3:0] p15 = (((5'd25)|(-3'sd1))*(-(-(2'd2))));
  localparam signed [4:0] p16 = {((-2'sd1)?(5'sd9):(2'd2)),{4{(3'd5)}}};
  localparam signed [5:0] p17 = (5'd21);

  assign y0 = (+{(&(~&((&p2)<<(!b3))))});
  assign y1 = (-(6'd2 * (a0>a0)));
  assign y2 = ($unsigned((($unsigned(b3))?$signed((-5'sd1)):(p6?a1:b3))));
  assign y3 = (+{{(-((~{p5,p17})<(p1<<<a5))),(-(-(!((+p16)|{p11}))))}});
  assign y4 = (2'd2);
  assign y5 = ((a2?b1:p2)?(b0?b5:a0):(5'sd11));
  assign y6 = ({b4,b4}<<(-(a2>p4)));
  assign y7 = (((-p2)>>(a3?a0:p9))>{{b4,p3}});
  assign y8 = (~(~|(-(a5&&b0))));
  assign y9 = (((b0===b3)?$signed(b5):{a5,b3})&$signed(((b3?a1:b4))));
  assign y10 = {4{p17}};
  assign y11 = (({b1,b5,b0}>>(-{{a3,b2,a5}}))===(|(6'd2 * (a1>=b1))));
  assign y12 = ((~^(!(~&(~^b0))))?((b3?p7:b1)?(~|p16):(b1?p3:a4)):(~&(p9?a0:b2)));
  assign y13 = (~^{p17});
  assign y14 = (-2'sd0);
  assign y15 = {3{((p15>>b4)&{4{p0}})}};
  assign y16 = (({3{p1}}?(p12<<<p9):{2{p6}})+((p16?b2:p14)<<<{4{a4}}));
  assign y17 = {2{(p16?a2:a5)}};
endmodule
