module expression_00483(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd3)<<(3'd7));
  localparam [4:0] p1 = (^(((2'd1)+(5'd17))>>((2'sd1)!=(4'd15))));
  localparam [5:0] p2 = (!(((4'sd3)<<(5'd23))>((3'd3)===(2'sd1))));
  localparam signed [3:0] p3 = ((3'd3)%(3'd4));
  localparam signed [4:0] p4 = (((4'sd4)?(4'sd1):(5'd23))?((+(2'sd0))^~((5'd6)?(3'sd1):(4'sd4))):((|(3'd0))==((5'd16)^(4'd10))));
  localparam signed [5:0] p5 = (({{(4'd9),(3'd6)}}<((5'd3)!==(3'sd1)))<=(((3'd0)<<<(-5'sd6))==((4'd12)!=(2'sd1))));
  localparam [3:0] p6 = ({3{(3'd5)}}|{4{(3'd1)}});
  localparam [4:0] p7 = (~|((!(+(~(|(5'd9)))))?(~&(~^(-((5'd29)*(2'sd0))))):(((3'd2)>(5'd9))>>>((3'd5)?(4'sd2):(3'sd1)))));
  localparam [5:0] p8 = (3'd4);
  localparam signed [3:0] p9 = (-((3'd7)?(-2'sd0):(-3'sd1)));
  localparam signed [4:0] p10 = (({(-4'sd4)}>>{3{(-2'sd0)}})+(5'sd12));
  localparam signed [5:0] p11 = (((2'd1)==(4'd10))&((4'sd3)!=(4'd13)));
  localparam [3:0] p12 = {3{(~&{4{(3'd3)}})}};
  localparam [4:0] p13 = (((+((-4'sd0)?(3'd4):(3'd2)))>(|((5'sd0)?(-2'sd1):(5'd27))))==(&((!(^(-5'sd8)))*((2'd0)?(5'sd4):(3'd6)))));
  localparam [5:0] p14 = {(^(-3'sd3)),((4'd0)&&(-3'sd0)),(6'd2 * (2'd2))};
  localparam signed [3:0] p15 = {2{{3{(-3'sd3)}}}};
  localparam signed [4:0] p16 = {1{(2'sd0)}};
  localparam signed [5:0] p17 = ((3'sd1)>>(2'd1));

  assign y0 = (4'sd6);
  assign y1 = ((~^{(a0|a1),(a5|a2),{b5,b3,a1}})?(~^((b2>b3)&{a3})):((b4||b4)<<<(~^{a2})));
  assign y2 = ((&(a1!==a4))||(b1|p3));
  assign y3 = ((^{3{b2}})>(~(&(!(a1^~b4)))));
  assign y4 = (b1&&b5);
  assign y5 = (6'd2 * (b0?b0:b2));
  assign y6 = ((a5&&b5)<(p7^~p8));
  assign y7 = ({(5'd7)}^~(4'd0));
  assign y8 = (-(!((~(~^(b1<<a2)))>((a5===a3)>>(~&b5)))));
  assign y9 = ((a2<<a0)!=(5'd27));
  assign y10 = (((4'd15)?(2'd1):(&a5))?$signed(((-(-a2))!={(&b5)})):(!(~|{{b0,b1,b2},(!p17),(^b0)})));
  assign y11 = (~((-b3)>>(b1<=a1)));
  assign y12 = (((b2===a2)?{1{p6}}:(p4>>>p12))?({(b2?a2:p2)}|{b2,p10,p12}):{3{(a3?a0:a2)}});
  assign y13 = (~&(^{{1{(!(!{{a2},(-b3)}))}},{2{{2{(~^p12)}}}}}));
  assign y14 = {1{{4{({4{b5}}>>(b3))}}}};
  assign y15 = {(~|{4{p8}}),{3{a5}},(p3^p17)};
  assign y16 = ((4'd13));
  assign y17 = (5'd2 * (p1<=p14));
endmodule
