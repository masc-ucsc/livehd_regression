module expression_00029(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(5'd28));
  localparam [4:0] p1 = ({1{(~^(((-3'sd0)!=(-4'sd3))<={(4'd12),(4'd12),(-3'sd3)}))}}!=={4{((3'd3)&&(4'd10))}});
  localparam [5:0] p2 = (|(+{(4'd13),(5'sd14)}));
  localparam signed [3:0] p3 = {4{(5'd17)}};
  localparam signed [4:0] p4 = {2{{{(3'd1),(2'sd0),(4'd0)}}}};
  localparam signed [5:0] p5 = {((-4'sd3)^~(5'd8)),((5'sd15)&(4'd9))};
  localparam [3:0] p6 = ((5'd9)-((2'd2)-(2'd3)));
  localparam [4:0] p7 = (|((5'sd1)&&(-5'sd1)));
  localparam [5:0] p8 = {1{(2'd0)}};
  localparam signed [3:0] p9 = (-2'sd1);
  localparam signed [4:0] p10 = (~&(|((((3'd7)&&(4'sd2))&(&(3'd6)))&&(3'd3))));
  localparam signed [5:0] p11 = {(&{(~(~{(2'sd1)})),(~{(2'd2),(2'd2),(-4'sd4)}),{(^(2'd0)),(~&(4'd6))}})};
  localparam [3:0] p12 = (4'sd5);
  localparam [4:0] p13 = (((~|(3'sd3))>((4'sd0)!=(-2'sd1)))||(~&(~(2'd2))));
  localparam [5:0] p14 = (4'd12);
  localparam signed [3:0] p15 = (3'd4);
  localparam signed [4:0] p16 = (((2'd2)^~(2'sd0))!=((3'd3)%(5'sd14)));
  localparam signed [5:0] p17 = ((!(^((-5'sd6)?(3'sd1):(3'd4))))?(-(!((3'sd3)?(-3'sd0):(5'sd4)))):(+((4'd1)?(5'sd2):(4'd11))));

  assign y0 = {((~$signed((p11)))<={a1,b0,p12}),($unsigned($unsigned((a3)))||((^p14)&&{p7,a4}))};
  assign y1 = ((~(!(&(~|p7))))^(!((2'd1)<(^b1))));
  assign y2 = ($unsigned({2{p3}})-(&{1{(p13?p4:p0)}}));
  assign y3 = ((!((^(p12+p16))<(a3!=a4)))|(({p10,p14,a5}||{1{p15}})==(b1?b3:a4)));
  assign y4 = {1{(3'sd0)}};
  assign y5 = {2{(b2?b3:b2)}};
  assign y6 = ((2'sd1)?(p12^b3):(b4==p7));
  assign y7 = {{{p9},{p5,b3}},{{a3,p12}}};
  assign y8 = {{4{p10}},{p16,p6,p3},(-(p8?p11:b1))};
  assign y9 = (p9^a2);
  assign y10 = (((b3>=a2)!=$signed(a1))?((b2?a1:b3)^~{b3,a2}):((b5)>=(a3<<<p9)));
  assign y11 = (((b4?b2:b5)?(a3?b5:p16):(3'd0))-(4'd13));
  assign y12 = (-3'sd0);
  assign y13 = ((&{p2,p16})==({p4,p10}>=(p3!=p4)));
  assign y14 = (((6'd2 * (6'd2 * p0))-($unsigned(p7)|{1{p3}}))^~((+(~&(~^a1)))===(~(b2^a5))));
  assign y15 = ({4{(~&b4)}}+{3{(~^{4{a1}})}});
  assign y16 = ((~|{p9,p12,p8})>={4{p0}});
  assign y17 = ((5'd2 * (p12?p0:p8))!=((p5!=p11)<(a3&&p8)));
endmodule
