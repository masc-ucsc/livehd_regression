module expression_00377(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd2)+(5'd2));
  localparam [4:0] p1 = {(-2'sd1)};
  localparam [5:0] p2 = (~&{{4{(2'd2)}},{(6'd2 * ((4'd2)>=(5'd21)))}});
  localparam signed [3:0] p3 = {(&{(5'sd0),(5'd16)})};
  localparam signed [4:0] p4 = ({1{((3'd7)<(4'd1))}}&(3'd3));
  localparam signed [5:0] p5 = (((5'sd12)?(-5'sd0):(4'd6))?(((3'd5)^(2'd2))||(5'd2 * (4'd7))):(((3'sd1)?(-4'sd7):(3'd5))-((5'd3)==(-3'sd3))));
  localparam [3:0] p6 = (!{{(2'd2),(-5'sd7),(-4'sd5)},{(-4'sd4),(2'sd0)},((5'd9)>=(5'sd9))});
  localparam [4:0] p7 = (!((((5'd19)>>(2'd0))?(&(3'd6)):((-5'sd9)?(5'd29):(-5'sd3)))<<(((4'sd2)>>>(3'sd1))?((-5'sd11)<<(3'd3)):((3'd0)?(2'sd0):(5'sd8)))));
  localparam [5:0] p8 = ((5'd2)<=(2'd0));
  localparam signed [3:0] p9 = ({2{(6'd2 * (4'd4))}}<<<(((-3'sd3)||(3'd4))?((-3'sd3)<<(5'd15)):((4'd11)?(-5'sd3):(2'd3))));
  localparam signed [4:0] p10 = ((((2'd2)+(2'd2))||((2'd0)?(4'd5):(-2'sd0)))<<<((+(3'sd1))||(5'd2 * (2'd3))));
  localparam signed [5:0] p11 = ((2'd2)?(-4'sd6):(-2'sd1));
  localparam [3:0] p12 = ({1{((4'sd2)==(3'd0))}}>>>(4'sd4));
  localparam [4:0] p13 = (({1{{1{((-3'sd0)<<(4'd14))}}}}&((4'sd4)>=((-3'sd3)===(-3'sd3))))===(((4'd4)>={4{(-2'sd1)}})<=(((4'sd3)==(5'd15))>((-3'sd0)|(-5'sd2)))));
  localparam [5:0] p14 = {((5'd9)<<<((5'd31)!==(2'sd1))),{{(4'd1)},((5'd30)&(5'd0)),(2'sd0)},(3'd3)};
  localparam signed [3:0] p15 = ((-4'sd1)^(((-3'sd3)&(4'd13))===((5'd25)?(5'd8):(-3'sd2))));
  localparam signed [4:0] p16 = ({1{((-5'sd7)<(2'sd1))}}?((4'd7)>(-2'sd1)):((4'd3)==(3'sd0)));
  localparam signed [5:0] p17 = (((-3'sd1)^(4'd11))-(^(~(3'd1))));

  assign y0 = {3{(&(-b5))}};
  assign y1 = ((b5?b2:a2)?((b1>=b2)|(a3?b2:a3)):$unsigned((a5!==b1)));
  assign y2 = {3{(({a4})<$signed({4{a5}}))}};
  assign y3 = {b3,p4};
  assign y4 = (~&((^({a4}))!==((b5!==b5)&(~|b2))));
  assign y5 = {3{(p8>p13)}};
  assign y6 = (5'd6);
  assign y7 = {(((p0?p14:a4))),{(|{a4,b3,p3})},{{(p14?p12:b0)}}};
  assign y8 = {3{(p16?a2:p10)}};
  assign y9 = (((b2?p8:p4)?(~|p5):$unsigned(p6))?{((p8)?(~&b4):(p1>>>p4))}:((b5!==a4)>>$unsigned((^p12))));
  assign y10 = {2{{3{p6}}}};
  assign y11 = (({3{{3{b2}}}}<=((5'd9)?(4'd13):{1{p16}}))<=(((3'd6)?(p6?a4:p3):{1{b1}})<<<(~(2'd0))));
  assign y12 = (~|((~&(&{2{a4}}))?(!(p8?b2:a2)):{p6,b3,a0}));
  assign y13 = (+{(!{1{{3{{p11,b1,b1}}}}})});
  assign y14 = (^(p13&b4));
  assign y15 = ((-2'sd0)>>(-(!(&(^(~&(^(3'sd1))))))));
  assign y16 = (!a5);
  assign y17 = (~^(+(|(~(((p11+p17)*(!a1))>>>(~(^(~|p8))))))));
endmodule
