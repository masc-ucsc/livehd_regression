module expression_00630(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {({(-3'sd3),(-5'sd11)}<<<{(4'sd0),(3'sd2)}),(((-4'sd3)?(5'd1):(2'sd1))<<((4'd9)?(5'd6):(-3'sd0)))};
  localparam [4:0] p1 = {{2{{1{{2{(-4'sd1)}}}}}}};
  localparam [5:0] p2 = (|(4'sd0));
  localparam signed [3:0] p3 = (((3'd2)?(-3'sd1):(4'sd1))?((-3'sd3)?(4'd4):(3'd2)):(2'd2));
  localparam signed [4:0] p4 = (((4'd10)-(3'sd1))^~(2'd0));
  localparam signed [5:0] p5 = {{{3{{4{(2'd0)}}}}}};
  localparam [3:0] p6 = ((((2'd3)&&(5'd28))>>>((3'sd1)===(2'sd1)))===(((2'd2)&(5'sd5))|((2'sd0)+(2'd0))));
  localparam [4:0] p7 = ((((3'd6)<=(-2'sd0))>>(|(-3'sd1)))?(2'sd1):(-3'sd2));
  localparam [5:0] p8 = (~(|(^(!(^(2'd1))))));
  localparam signed [3:0] p9 = (~|((((5'd29)?(-2'sd0):(-5'sd8))==((2'd3)>(3'd4)))==(((4'sd3)^(5'd18))+((5'd3)?(-3'sd2):(3'sd3)))));
  localparam signed [4:0] p10 = (((-5'sd9)?(2'sd0):(4'd7))?{(3'd0)}:((3'sd3)+(-2'sd1)));
  localparam signed [5:0] p11 = ((~&{3{(5'sd2)}})-(~^{2{(2'd3)}}));
  localparam [3:0] p12 = {(~|((3'd2)^(5'd5))),(~(!(-(-2'sd1)))),(|(~&((3'd4)-(2'd2))))};
  localparam [4:0] p13 = {3{((-5'sd11)?(2'd0):(3'd2))}};
  localparam [5:0] p14 = (&((-(|(5'd2 * (3'd3))))>>(~&(-3'sd0))));
  localparam signed [3:0] p15 = (~^((((-5'sd1)+(3'd7))<=((2'sd0)!=(4'd8)))>=((~^(-(-5'sd7)))<=((2'd3)&(-5'sd0)))));
  localparam signed [4:0] p16 = ((((5'd18)<=(3'd6))>((-2'sd0)<=(2'sd1)))<<(-({(-3'sd2),(-5'sd7),(2'd2)}>>>((3'sd3)^(2'sd1)))));
  localparam signed [5:0] p17 = (4'd2 * ((2'd2)||(3'd1)));

  assign y0 = (&{(~&(~|(~(~(p16?b1:p11)))))});
  assign y1 = (~&((!(b0==p4))^~((p1>p8)+(p7>>p14))));
  assign y2 = (|(~|{4{(&p4)}}));
  assign y3 = (((2'd2)&&(|(2'd1)))?((a3>>p7)?{b1,b5,b2}:(~&a0)):((a5?a5:b2)<<{{3{b5}}}));
  assign y4 = ($unsigned((+((~^{$signed(b4)})^~((4'sd0)<<<(p11)))))-{{a0,b0,b5},(a5^~p16),(4'sd0)});
  assign y5 = $signed($unsigned((($signed((b0?p0:p15))>>>$signed({b4}))||((b5?p4:p0)?{p15,p17,b3}:(p8<<p11)))));
  assign y6 = (|(((4'd9)?(p6||a1):(|p11))?($signed((p1&&p15))<=$unsigned((p9))):$unsigned((-3'sd3))));
  assign y7 = {3{p13}};
  assign y8 = (3'd6);
  assign y9 = ((p10?b1:a4)?{4{p15}}:(p9?p10:p5));
  assign y10 = (|(3'sd1));
  assign y11 = {4{p1}};
  assign y12 = (((p12>>p3)+(+(p14>p11)))+(+{4{b0}}));
  assign y13 = ((~|$unsigned((|b0)))>>>((^$signed(b5))));
  assign y14 = (((p11&p8)<=(p10<p3))>=((p5&p8)>(p4-p8)));
  assign y15 = ((a3===a3)&(a4!=p6));
  assign y16 = ($unsigned((((a0!==a0)||$unsigned(b2))^((a4)|(p13==p16))))||$unsigned(((2'd2)&&(3'd6))));
  assign y17 = ((-3'sd0)!=(-4'sd7));
endmodule
