module expression_00310(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(((~|(-4'sd2))!=((2'sd0)>>>(5'd1)))>>>(((-4'sd1)>>>(-4'sd7))^~((3'sd2)<<<(2'd1)))));
  localparam [4:0] p1 = (&((2'd3)|(!{((3'd4)-(5'd17)),{(4'sd7),(-2'sd0)}})));
  localparam [5:0] p2 = ((((-5'sd5)>(-2'sd0))&&((-4'sd3)<<(5'd12)))?(&((2'd2)?(-2'sd1):(5'd0))):{((|(-4'sd6))&&{(-4'sd3),(-2'sd0)})});
  localparam signed [3:0] p3 = (2'd3);
  localparam signed [4:0] p4 = (((3'sd0)-(5'd16))!==((3'sd2)>=(3'd2)));
  localparam signed [5:0] p5 = {{((5'd28)&(-2'sd0))},((-2'sd0)?(2'd3):(5'sd1)),({(3'sd1)}&{(2'sd1),(3'sd1)})};
  localparam [3:0] p6 = (((-3'sd3)?(2'd0):(-5'sd11))?{(-2'sd1),(2'd0),(-4'sd2)}:((-2'sd0)>>>(5'd23)));
  localparam [4:0] p7 = ((-3'sd0)>>(-5'sd3));
  localparam [5:0] p8 = (|((((2'd3)>>>(4'd14))%(-2'sd1))||((~^((-4'sd2)-(-2'sd1)))>(&((2'sd0)^~(-2'sd0))))));
  localparam signed [3:0] p9 = ((2'sd1)<<(3'sd0));
  localparam signed [4:0] p10 = (^((~(~|((-5'sd5)>(-3'sd3))))||(&(((3'd3)>=(4'd1))===((3'd4)<=(3'sd0))))));
  localparam signed [5:0] p11 = (~^(-2'sd0));
  localparam [3:0] p12 = ((2'sd1)?(4'd1):(5'd16));
  localparam [4:0] p13 = ((2'd1)<<<(2'd1));
  localparam [5:0] p14 = {((4'd9)?(-5'sd13):(2'd1)),((2'd1)?(-3'sd0):(2'd2)),(~|((-5'sd15)===(2'd2)))};
  localparam signed [3:0] p15 = (~{1{({1{(+((^(5'd22))>(&(-4'sd4))))}}^~{2{{1{(^(5'd9))}}}})}});
  localparam signed [4:0] p16 = ((3'd2)|(2'sd1));
  localparam signed [5:0] p17 = (+(((+(-2'sd1))>>>(5'sd11))+(5'd25)));

  assign y0 = (a5?a1:b2);
  assign y1 = (((p10?p15:p9)^~(b4?p7:b1)));
  assign y2 = ($signed(((b3?p9:a4)))?($signed(b3)?$signed(p4):(b1)):$unsigned(((p0?a2:b5))));
  assign y3 = ((6'd2 * (6'd2 * p2))<(~^(+(4'd2 * (2'd2)))));
  assign y4 = {3{{1{((p6||p1)&{1{p5}})}}}};
  assign y5 = (5'sd10);
  assign y6 = ((5'd26));
  assign y7 = {4{(a0?b0:b4)}};
  assign y8 = {3{{2{(p14|p3)}}}};
  assign y9 = {1{((-3'sd2)<=(p5!=p1))}};
  assign y10 = (~&(5'd2 * (~^$unsigned(a2))));
  assign y11 = ((~^p15)?(~^p3):(&a4));
  assign y12 = (((b4>>p17)?(p15>>>a1):(a2>>p11))?((p17?p4:a2)-{3{p0}}):((~&(p11?p13:p11))<=(p8?p4:p4)));
  assign y13 = (~&(-2'sd0));
  assign y14 = {(2'sd0),{4{b1}},$signed((p10>p3))};
  assign y15 = {({p16,b4}<=(p16>=a3)),{{(b2>=b1)}},((~^b1)!=={a4})};
  assign y16 = ({(p17?p17:p12),(4'd3)}?(-2'sd1):(3'sd0));
  assign y17 = ($unsigned((-3'sd3))!={p12,p15,p7});
endmodule
