module expression_00117(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({2{(2'sd1)}}?((-2'sd1)+(-4'sd2)):((-4'sd2)?(5'sd7):(3'sd2)))>>({3{(-5'sd1)}}<=((3'sd0)^~(-5'sd2))));
  localparam [4:0] p1 = (((5'd18)&(5'd10))?(5'd2 * (4'd1)):((3'sd1)||(4'd3)));
  localparam [5:0] p2 = (|(((2'd0)?(5'd12):(4'sd7))?(5'd26):((-5'sd3)?(2'd1):(3'd1))));
  localparam signed [3:0] p3 = (((5'sd5)>=(2'sd1))||((-2'sd0)&&(3'd1)));
  localparam signed [4:0] p4 = {((2'd3)&(-5'sd1))};
  localparam signed [5:0] p5 = (-(^(!(~|(+(~(-3'sd2)))))));
  localparam [3:0] p6 = {(4'sd7)};
  localparam [4:0] p7 = (6'd2 * ((2'd1)^~(5'd19)));
  localparam [5:0] p8 = (((&((4'sd6)?(-3'sd3):(-2'sd1)))<(~^(~(4'd15))))>>(!(4'd3)));
  localparam signed [3:0] p9 = (((4'd11)-(-3'sd0))*(~&(^(4'd7))));
  localparam signed [4:0] p10 = {(-4'sd0),(4'sd2)};
  localparam signed [5:0] p11 = {{{3{((3'sd2)-(5'd27))}}}};
  localparam [3:0] p12 = {((-3'sd3)<<(3'sd2)),{(-5'sd8),(3'd6),(4'sd6)}};
  localparam [4:0] p13 = ((((2'd0)===(3'sd3))<((4'd4)<<(5'sd6)))|(3'd6));
  localparam [5:0] p14 = ((!(5'd23))>={3{(5'd24)}});
  localparam signed [3:0] p15 = (-((+(2'd2))&&({(3'sd0)}==((2'd1)<<(2'd0)))));
  localparam signed [4:0] p16 = ({{(-3'sd1),(2'sd0)}}?(^(+(~^(2'sd0)))):(~&((2'd3)>=(3'd0))));
  localparam signed [5:0] p17 = ((3'd2)?(3'd3):(3'sd1));

  assign y0 = (({{(a3-b0)},(6'd2 * p1),(a4!=b1)})>((~&(a0!=p8))>$unsigned((a3>>>p12))));
  assign y1 = $signed({p7,p5,p10});
  assign y2 = (~&({1{{3{{4{b5}}}}}}^~((|{4{p3}})^~(~|(~|b2)))));
  assign y3 = (((b3^b1)!==(6'd2 * b2))&&{(6'd2 * b2),{4{b0}},(b0<<a3)});
  assign y4 = ((-{3{{3{a2}}}})+{2{({p14}<={2{p6}})}});
  assign y5 = (((-((&b1)?$unsigned(a2):(a0?a3:b5)))?($signed(b4)?(-2'sd1):(5'd9)):(+(2'd2))));
  assign y6 = (-5'sd8);
  assign y7 = ({{4{b3}},(^(^p2)),{p15,p16}}&&{2{(&{1{(p7>>>p10)}})}});
  assign y8 = (6'd2 * (p7?p8:p14));
  assign y9 = (((p4<<<p16)?(p9?p1:p13):(p8?p15:p14))<$unsigned(((p10||p10)?(4'sd6):(2'd2))));
  assign y10 = {3{{3{(b0>>>b1)}}}};
  assign y11 = (((~&a0)^(a4!=a3))^{b5,b0,b5});
  assign y12 = {4{(^(^(-3'sd0)))}};
  assign y13 = ((!{(a4!==a1),{a5,a3,a5}})<<{({(-5'sd3)}<<<(5'sd3))});
  assign y14 = $signed({3{(~^(p14?a1:p12))}});
  assign y15 = (p5?p4:p1);
  assign y16 = (+(&(~|(~|((5'sd8)!=((a3+a3)=={2{p17}}))))));
  assign y17 = (&$signed((2'd3)));
endmodule
