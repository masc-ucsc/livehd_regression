module expression_00986(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{3{(((4'd4)>(5'd7))&&(|(4'd1)))}});
  localparam [4:0] p1 = (!(-5'sd14));
  localparam [5:0] p2 = {2{{2{{{(3'd1)}}}}}};
  localparam signed [3:0] p3 = (!(+(&((-(-5'sd12))>>(-5'sd10)))));
  localparam signed [4:0] p4 = (((4'd9)>>(3'd2))>>((-4'sd5)!==(5'd10)));
  localparam signed [5:0] p5 = {3{((-3'sd2)<(-5'sd9))}};
  localparam [3:0] p6 = ({1{((3'sd2)<(5'd22))}}<<{3{(5'd22)}});
  localparam [4:0] p7 = ((-2'sd0)|(3'sd2));
  localparam [5:0] p8 = (-3'sd3);
  localparam signed [3:0] p9 = (~^{(((3'sd1)<<<(4'd12))==(!(5'd21)))});
  localparam signed [4:0] p10 = {2{(!{2{{{(4'd11)}}}})}};
  localparam signed [5:0] p11 = {({{(((2'd2)==(-5'sd2))&&((4'd3)===(-5'sd10)))}}>>>(((-4'sd7)+(2'sd1))^((-4'sd4)!==(3'd3))))};
  localparam [3:0] p12 = (~(2'd2));
  localparam [4:0] p13 = ((5'd6)!=(4'sd5));
  localparam [5:0] p14 = (-(~^(((4'sd6)<=(3'd4))>>>((3'd0)<(3'sd0)))));
  localparam signed [3:0] p15 = {{3{(4'd6)}},(~|{3{(-3'sd0)}})};
  localparam signed [4:0] p16 = (((~&(-3'sd2))!=((4'd3)?(-3'sd0):(3'd1)))?((5'sd8)===(!(3'sd2))):((5'd10)?(-5'sd14):(-4'sd3)));
  localparam signed [5:0] p17 = (2'd3);

  assign y0 = ((&(((^p1)<<(p5|p5))<=(6'd2 * (~^p1))))+(+(({p14,p11}>>(p16^~p15))<(|(p0^p8)))));
  assign y1 = ((4'd2 * (p14<<p1))<((b0!=a1)!==(b3<b2)));
  assign y2 = (~&(5'd1));
  assign y3 = (4'd5);
  assign y4 = (((a4?a1:b2)?(p8<a4):(+(p17-b4)))>=(!((b2<=b0)?(~|p2):(&p3))));
  assign y5 = ({1{$signed((b5-b5))}}<<((p8|b5)>{4{b4}}));
  assign y6 = (((b3?p0:a1)?(~&(p16%p6)):(|(p16-b4)))<<<(((a0||b3)!==(a2<<b2))<<((b2&&p6)>>(p3?b4:a4))));
  assign y7 = ((a2-b0)!==(4'd5));
  assign y8 = (-2'sd0);
  assign y9 = (~^({3{a2}}?$signed((^(p3?p10:p15))):(p6?p7:p0)));
  assign y10 = $signed(({a0,a5,a0}?{a3,b4}:(4'd13)));
  assign y11 = (4'sd5);
  assign y12 = $signed(((b3?b4:a0)?(b3?b4:b3):(b4?a1:a0)));
  assign y13 = {3{({1{b0}}>(p9|b4))}};
  assign y14 = (((p12+p14)+(b4>>b4))<{4{(a4+p7)}});
  assign y15 = (5'd26);
  assign y16 = (((p2?p11:p13)?(p3||p1):(p17^~p13))&($signed($unsigned(p12))?(p0<<p10):(p1?p15:p5)));
  assign y17 = $signed(p15);
endmodule
