module expression_00096(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&((5'd18)<(-4'sd0)));
  localparam [4:0] p1 = (((3'd1)<<(3'd3))||((2'd3)||(5'd15)));
  localparam [5:0] p2 = ((~^((5'sd5)^(5'd22)))|{(!(2'd2))});
  localparam signed [3:0] p3 = (!((((5'd3)>(4'd14))<<(|(5'd10)))!==(~(6'd2 * (5'd26)))));
  localparam signed [4:0] p4 = (~&(-4'sd7));
  localparam signed [5:0] p5 = (((5'sd11)>>(5'sd9))||(-(2'd3)));
  localparam [3:0] p6 = ((3'd5)?(((4'd5)>>>(5'd0))-((2'd3)!==(5'd8))):((5'd26)===(~&(-2'sd0))));
  localparam [4:0] p7 = (((((3'sd2)>(-2'sd0))<(~^(4'd2)))<(~((5'sd5)<(3'd1))))<<((~^((3'sd2)===(3'd1)))==(!((4'sd0)-(3'sd2)))));
  localparam [5:0] p8 = {{(4'sd3),(5'd26)},(~|(5'd31)),((2'd3)?(5'd4):(-2'sd0))};
  localparam signed [3:0] p9 = {(|(5'd2 * {(4'd2 * (4'd3))})),({1{(-4'sd1)}}?(6'd2 * (5'd6)):((4'd15)?(4'sd7):(-5'sd2)))};
  localparam signed [4:0] p10 = (4'd15);
  localparam signed [5:0] p11 = ((3'sd0)-(2'd0));
  localparam [3:0] p12 = (+(|(((3'd7)+(2'sd0))!==((5'sd10)==(4'd11)))));
  localparam [4:0] p13 = ((~|((3'd3)?(-4'sd7):(4'd3)))?{1{{3{(-5'sd11)}}}}:{2{(+(-3'sd2))}});
  localparam [5:0] p14 = (!(&(-(^(-3'sd0)))));
  localparam signed [3:0] p15 = ((2'sd1)-(5'sd1));
  localparam signed [4:0] p16 = (5'd2 * {1{((2'd3)<<<(5'd30))}});
  localparam signed [5:0] p17 = {4{(((3'd2)<(4'd4))^{4{(4'd6)}})}};

  assign y0 = {a1};
  assign y1 = (p5||a5);
  assign y2 = (&{2{((~p1)>>>$unsigned(b1))}});
  assign y3 = (~^(-4'sd7));
  assign y4 = {{3{a3}},(5'd2 * $unsigned(a2)),{a5,a2,a3}};
  assign y5 = (3'd4);
  assign y6 = ({4{b2}}&(a3<a3));
  assign y7 = ({1{(a5!==b0)}}?(~|(b4?p7:p4)):(~(3'sd3)));
  assign y8 = ((~b5)^(b2|b2));
  assign y9 = (~^(~^{(b5>>b5),(a0<<<a2),(-p11)}));
  assign y10 = (|(({(5'sd2),(|a4)}&&((2'sd1)||{1{a2}}))-{(^{(b4?b3:a4),$signed(a1),(a3<b1)})}));
  assign y11 = {(p15?p10:p13)};
  assign y12 = ((~|$unsigned((((($unsigned((p1<=b4))))))))<=($signed((^(^(a1<b4))))===((~a2)<=(b2<<<b4))));
  assign y13 = ((p13?p2:p10)?(p3==p7):(|p11));
  assign y14 = ((&(3'd2))^~((b5^~a1)=={1{p11}}));
  assign y15 = (-$signed({((!(-$signed((({b4,a1}||(&a1))))))<{(~(-(~|(~(&(&(b5|a2)))))))})}));
  assign y16 = (((a2%p6)<<(a0?b1:p9))||(&((~|p4)?(~p3):(|p0))));
  assign y17 = (((p7+p16)^~(p5||p8))^~(4'sd4));
endmodule
