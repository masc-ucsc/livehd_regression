module expression_00034(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-3'sd3)==(-(-4'sd4)));
  localparam [4:0] p1 = ({((5'd22)||(3'sd0)),((5'sd1)^~(5'd3)),((3'sd1)?(-3'sd2):(-5'sd11))}&(((4'd12)?(3'd1):(4'd12))?{(3'sd0)}:((4'd0)>(-4'sd1))));
  localparam [5:0] p2 = (+{(&(2'd1)),{(4'sd4)}});
  localparam signed [3:0] p3 = (4'd1);
  localparam signed [4:0] p4 = {(&{{1{{(4'd9),(5'd27)}}},(!(&(!(5'd25))))})};
  localparam signed [5:0] p5 = {{((-2'sd1)^(-2'sd1)),(|(3'd2))}};
  localparam [3:0] p6 = ((((5'sd0)===(3'd1))>=(-(-2'sd0)))<=((~&(4'd3))||(-4'sd6)));
  localparam [4:0] p7 = {((-5'sd0)?(-3'sd0):(4'd3)),{(2'd1),(-3'sd2)}};
  localparam [5:0] p8 = {4{(-4'sd3)}};
  localparam signed [3:0] p9 = {(^{4{((4'd8)^(4'd5))}})};
  localparam signed [4:0] p10 = (((2'sd0)?(3'sd1):(5'sd15))?{1{(3'sd3)}}:{2{(4'd2)}});
  localparam signed [5:0] p11 = (-5'sd6);
  localparam [3:0] p12 = {((3'd6)?(4'd14):(2'sd0)),{(5'sd0)}};
  localparam [4:0] p13 = {4{(2'd1)}};
  localparam [5:0] p14 = ((~(3'd5))?((-3'sd2)!==(-4'sd7)):((2'd0)?(-5'sd1):(2'd2)));
  localparam signed [3:0] p15 = (((4'd15)?(5'sd0):(3'd5))?((4'd14)?(2'd1):(2'd0)):((2'sd0)?(4'd8):(4'd3)));
  localparam signed [4:0] p16 = ({((3'd5)===(4'd9)),(2'd2),(5'd2 * (4'd9))}>{(-(3'd7)),(2'd3),(&(2'sd1))});
  localparam signed [5:0] p17 = {1{((!(~^(-(^(2'sd1)))))?{4{(4'sd1)}}:{3{(~&(5'sd11))}})}};

  assign y0 = ((p11^p17)?(a0!==a2):(b3|p11));
  assign y1 = (~(({p8,p6,p11})-{(p0==p16)}));
  assign y2 = (5'd2 * (a2<<<a2));
  assign y3 = (-({3{(p15?b0:p5)}}||((b3&b2)?(b5&p1):(a3&p1))));
  assign y4 = (3'sd0);
  assign y5 = (((~|p15)?{p4,p9,p11}:(~&p14))?{(&p14),(p12<p6),(|p10)}:(4'd2 * (p14>>p13)));
  assign y6 = (!($signed((5'sd9))?(~(5'd31)):{{2{p6}}}));
  assign y7 = {(p0<<<a3)};
  assign y8 = (((-2'sd0)==(p1>=p11))<((2'sd1)-(5'd11)));
  assign y9 = $unsigned($signed((~^(a2))));
  assign y10 = (&(~|(~|(~^p2))));
  assign y11 = (((b3?p6:a4)?(|p6):(~|p12))?(-(^$signed((p16?a3:p17)))):(!(|$signed({{p7,b0},(p6<=p3)}))));
  assign y12 = (-3'sd0);
  assign y13 = $unsigned(((a1-a0)===$signed($unsigned(a3))));
  assign y14 = ((4'd2 * (a1>>>a0))!==(((b0!=b5)<(a0>=b3))>=((a3<<<b4)<<(b3==a3))));
  assign y15 = (~^(b1?p4:p5));
  assign y16 = (((-(b4!==b0))<<{2{(a4>=p15)}})^((~&(-3'sd1))-((&p7)&&(p17>>>p9))));
  assign y17 = (2'sd0);
endmodule
