module expression_00824(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(({4{(-3'sd3)}}?((5'd7)?(4'd6):(4'sd2)):{2{(3'd3)}})?{3{{(4'd5)}}}:({4{(4'd7)}}?{(4'sd3)}:{(-4'sd2),(-4'sd0),(-5'sd5)}))};
  localparam [4:0] p1 = ({(2'sd0),((4'd1)+(2'd1))}?(((3'sd1)?(3'sd0):(-3'sd2))?{(2'd1)}:(~(5'sd6))):(((5'd18)<(-5'sd11))||(5'd10)));
  localparam [5:0] p2 = {{{(4'd0),(2'd3),(3'd5)},(~|{(4'd6),(4'sd6)})}};
  localparam signed [3:0] p3 = ((5'd20)>>>(5'd0));
  localparam signed [4:0] p4 = {3{((5'sd1)?(3'd3):(-4'sd2))}};
  localparam signed [5:0] p5 = ((3'd2)<<<(4'd10));
  localparam [3:0] p6 = ({4{(-3'sd1)}}?((4'sd1)>>(-3'sd2)):{1{{(-5'sd8)}}});
  localparam [4:0] p7 = (-{(+(((|(~&(-2'sd0)))&&(-{4{(3'd2)}}))|(!(-4'sd1))))});
  localparam [5:0] p8 = {2{(-5'sd2)}};
  localparam signed [3:0] p9 = ((3'd6)?((3'd4)?(-5'sd11):(4'sd3)):(~(~&(~(4'd15)))));
  localparam signed [4:0] p10 = (&(~|{(|((-5'sd3)!=(5'd8)))}));
  localparam signed [5:0] p11 = ((~|(~|((-2'sd0)!==(4'sd7))))>>(~(|(~|(3'd2)))));
  localparam [3:0] p12 = ((&(4'd15))!={4{(4'd1)}});
  localparam [4:0] p13 = {{(2'd1),(5'd5),(5'd14)},(3'd7),((5'd27)>(3'd4))};
  localparam [5:0] p14 = (|((((3'sd3)-(4'sd2))<((2'd3)>=(4'd6)))=={((2'd0)?(4'd3):(5'd7)),{(-3'sd3)},((5'd28)&&(3'd6))}));
  localparam signed [3:0] p15 = (^{3{(2'sd1)}});
  localparam signed [4:0] p16 = (4'd2 * ((2'd3)?(3'd6):(4'd7)));
  localparam signed [5:0] p17 = {4{(!{1{{1{(2'd0)}}}})}};

  assign y0 = {{((b3&a4)>>>(a5<a2)),(4'd2 * (a1^~a2)),({b5,b4,b5}&&(a5<<b4))}};
  assign y1 = ((~&{3{(&b2)}}));
  assign y2 = ((2'sd1)&(((|b1)===(a0>>a4))>((~&p1)>>(~|p13))));
  assign y3 = (3'd3);
  assign y4 = ($signed((a0?p12:a5))||(^(a0>>a2)));
  assign y5 = ((p10&&p2)?$unsigned(a0):(p17%p1));
  assign y6 = (((4'sd3)&&(p11^b2))!=(-4'sd3));
  assign y7 = {$unsigned((!((p15?p7:p16)?(b2):(~&p11)))),((~|(p2))?(p4?p8:a0):((~|p12)))};
  assign y8 = (4'd2 * {4{b0}});
  assign y9 = $signed((|(({1{$unsigned(a0)}}<=(~$unsigned(a5)))>>>$signed(((p9>b0)<<<(~&(p13)))))));
  assign y10 = (~|{4{(~^{4{p5}})}});
  assign y11 = {1{{3{{(b0?p1:p14),{2{a1}},{1{b5}}}}}}};
  assign y12 = (!(((p10<b1)<(b1!==b5))<=$unsigned((-(a4>p8)))));
  assign y13 = ({2{(((p9?b2:b1)?(b1?p10:b2):(~^p2)))}});
  assign y14 = {$unsigned((&(((~^p11)<(a4!==b5))<={(-p16),{p6}}))),(((p1<p1)>>>{p2})+((b5>a5)+(p10>>p14)))};
  assign y15 = (-3'sd3);
  assign y16 = $unsigned((+$signed($unsigned((+((b1===b4)))))));
  assign y17 = (({3{p2}}?(b1-b2):{a5})?((b1&&p1)>={b5,a3,a5}):{((p9?b3:b2)?(4'd2 * a0):(b1?b2:b0))});
endmodule
