module expression_00005(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(&(!(-(&(!(&(-4'sd0))))))));
  localparam [4:0] p1 = (((5'd27)==(-3'sd0))/(5'sd8));
  localparam [5:0] p2 = ({1{{4{(3'sd1)}}}}<{4{(4'd13)}});
  localparam signed [3:0] p3 = {{2{(2'sd0)}},{3{(5'sd9)}},{{(3'd6)}}};
  localparam signed [4:0] p4 = {((((3'sd1)>>(5'd3))<=((5'd8)+(2'sd1)))^{(4'd8),(-4'sd6),(3'sd2)})};
  localparam signed [5:0] p5 = (^{1{(~|(~{2{{1{(~{2{(4'sd5)}})}}}}))}});
  localparam [3:0] p6 = (^(&(4'd0)));
  localparam [4:0] p7 = {3{((4'd6)&(3'sd3))}};
  localparam [5:0] p8 = ((((5'sd13)|(2'd0))>((3'd6)^~(3'sd1)))==({(5'd15),(2'd1),(2'd2)}&&((-2'sd1)>(5'd15))));
  localparam signed [3:0] p9 = ((-5'sd12)<<(5'd0));
  localparam signed [4:0] p10 = (3'd2);
  localparam signed [5:0] p11 = (((6'd2 * (3'd4))?((5'd21)<=(-4'sd1)):((2'd3)+(4'sd4)))?(~((^(5'd24))>=(|(4'd12)))):(((3'sd0)-(2'd1))^~((4'd6)?(3'd0):(4'd7))));
  localparam [3:0] p12 = (|(6'd2 * ((3'd2)?(3'd4):(3'd4))));
  localparam [4:0] p13 = ((&((-3'sd1)>>(-3'sd3)))^((!(2'd0))^((-4'sd5)<<(4'sd0))));
  localparam [5:0] p14 = (((4'sd0)?(4'd6):(2'sd0))<({1{(-2'sd0)}}>>>{4{(2'd3)}}));
  localparam signed [3:0] p15 = (((3'd0)!==(3'sd3))<((5'd20)?(5'd9):(-2'sd0)));
  localparam signed [4:0] p16 = (({1{(-4'sd5)}}>(~|(4'sd0)))<({4{(2'd2)}}<((-5'sd1)<=(3'sd3))));
  localparam signed [5:0] p17 = (|(~(4'sd3)));

  assign y0 = $unsigned({3{({3{p16}}<=$unsigned(p17))}});
  assign y1 = {2{{{(4'sd4),(3'd3),{2{a4}}}}}};
  assign y2 = (-(~^(!{{{2{b3}},{4{p5}}}})));
  assign y3 = (+(&(|(!(+(-(5'sd2)))))));
  assign y4 = (|(|(b4?a0:a3)));
  assign y5 = ((3'sd3)<(2'd1));
  assign y6 = ((+(&({1{a2}}<<<{4{p4}})))^~((5'd4)>>{4{p3}}));
  assign y7 = {3{b1}};
  assign y8 = {3{{2{a5}}}};
  assign y9 = (~&(|(~(+(-(+(&(|(!(^(~&(^(-(&(~(~(&(+(!(~&p0))))))))))))))))))));
  assign y10 = (((p3==p15)<={a2,a1,a3})>=(~&(~^{b1,p16,b4})));
  assign y11 = (~&(2'd0));
  assign y12 = (3'd3);
  assign y13 = ((!{2{(p0?p9:a5)}})?((p2^b3)<={1{(a4>>>p10)}}):((b5^~p4)>(a3!=b3)));
  assign y14 = ({{b2,a3,b3},(a2?a1:a1),(a5&&a2)}>={{(a0?b1:b0)},(~|((a1?a5:b1)!=(b0?b5:b5)))});
  assign y15 = (^a5);
  assign y16 = (~^(-b1));
  assign y17 = (a2?p6:p7);
endmodule
