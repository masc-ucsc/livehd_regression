module expression_00528(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+((3'sd2)&&(2'sd0)))?(^(4'd5)):((-4'sd3)?(-4'sd4):(5'd2)));
  localparam [4:0] p1 = (!({((2'sd1)!==(4'd1)),((2'd3)+(-4'sd6))}^{(-2'sd1),(5'd9),(2'sd1)}));
  localparam [5:0] p2 = (~^{1{{3{(~&(3'd7))}}}});
  localparam signed [3:0] p3 = ((&((2'd3)?(5'd10):(5'd18)))?{4{(-3'sd2)}}:{1{(^(-3'sd0))}});
  localparam signed [4:0] p4 = ((4'd5)?(3'd1):(2'd0));
  localparam signed [5:0] p5 = (|{(^(-5'sd3)),(~|(5'd29)),(~|(4'd10))});
  localparam [3:0] p6 = ((((4'sd6)<=(4'd4))<<((2'd3)|(4'd15)))?(((-5'sd1)<(-5'sd11))?{(3'd5),(2'd1)}:((5'sd6)!=(4'd6))):(((5'd9)===(-5'sd11))?((-5'sd3)<<(-2'sd1)):((4'd11)<<<(2'd3))));
  localparam [4:0] p7 = {1{{4{((4'sd1)^(-4'sd3))}}}};
  localparam [5:0] p8 = {1{(((4'd4)&&(-3'sd0))?(4'd2 * (3'd0)):((-5'sd0)?(3'd6):(3'sd3)))}};
  localparam signed [3:0] p9 = ((((2'sd1)===(4'sd2))%(4'd8))!=(4'd2 * ((2'd0)&&(2'd3))));
  localparam signed [4:0] p10 = {1{(^(4'd8))}};
  localparam signed [5:0] p11 = ((-((3'sd2)<<<(3'd0)))*(4'd7));
  localparam [3:0] p12 = {3{(2'd0)}};
  localparam [4:0] p13 = {(((4'd12)===(2'sd0))&((3'd4)<(4'sd5))),{({(5'd15),(-2'sd0)}>>>((2'sd1)>>>(3'sd0)))}};
  localparam [5:0] p14 = ({3{(2'd1)}}|{4{(2'd1)}});
  localparam signed [3:0] p15 = ((6'd2 * (2'd2))?((-5'sd4)<=(4'sd6)):(+{(3'sd3),(-3'sd2),(3'd5)}));
  localparam signed [4:0] p16 = (-5'sd12);
  localparam signed [5:0] p17 = ((-(((5'd13)>=(5'd22))&((2'd2)<=(3'd7))))<=(((3'd5)!=(3'd2))!==((5'sd11)<(4'd12))));

  assign y0 = (!(~&($unsigned(p16)>>(b2-a4))));
  assign y1 = (((p16?p7:p10)&&(p3?p16:p17))<<(+(|(4'd2 * p13))));
  assign y2 = (3'sd1);
  assign y3 = (3'd3);
  assign y4 = (~|{({p16,p15,p2}?(^p8):{b3,p15}),{3{(p7<=p10)}}});
  assign y5 = (5'd1);
  assign y6 = {(-{{3{p7}},(a1===b1),(a3&&p11)})};
  assign y7 = $unsigned($signed({3{$signed((~p5))}}));
  assign y8 = {3{b0}};
  assign y9 = (5'd2 * (!(p8>>p8)));
  assign y10 = {{4{{b1,a3}}},(!{(!(a2>>b5))}),((b0===b2)<=(~|(b4&&a4)))};
  assign y11 = {4{{4{p11}}}};
  assign y12 = {2{b1}};
  assign y13 = {((p10<p1)^(a0>>>a3)),{4{(a4===a1)}},(-5'sd4)};
  assign y14 = {2{(2'd2)}};
  assign y15 = (|(4'sd4));
  assign y16 = (4'd11);
  assign y17 = ((b3==a4)?(a0?a3:a1):(p0<<<a4));
endmodule
