module expression_00239(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((|((5'sd11)>>(4'd0)))||((-5'sd15)!==(3'd6)));
  localparam [4:0] p1 = (-{{(4'd9)},(~|(2'd3)),((3'd1)?(2'sd1):(5'sd6))});
  localparam [5:0] p2 = ((+(~^(4'sd2)))?(~|((3'sd2)&(3'd6))):(-(~|(-3'sd2))));
  localparam signed [3:0] p3 = ((|((~|(2'd3))==={2{(-3'sd2)}}))^(~|(((5'd24)|(3'd7))!=((-4'sd6)>>(3'd3)))));
  localparam signed [4:0] p4 = ((((-4'sd5)%(2'd1))||((4'd11)%(-4'sd2)))>=(~|((|(-2'sd1))>=(!(5'd12)))));
  localparam signed [5:0] p5 = (((~((-4'sd0)?(2'd1):(3'sd0)))>((-3'sd2)>>>(-4'sd3)))>>(((4'sd3)?(-5'sd13):(2'sd1))|((4'd7)<=(5'd21))));
  localparam [3:0] p6 = {{(((3'sd3)===(2'd3))-{(3'd6),(-4'sd0),(5'd9)}),(((-5'sd2)<<<(4'sd1))^~((5'd16)!==(-3'sd3))),{3{(-4'sd6)}}}};
  localparam [4:0] p7 = {3{(-2'sd0)}};
  localparam [5:0] p8 = {{{3{{4{(2'd0)}}}}}};
  localparam signed [3:0] p9 = {4{{(3'd1),(3'd0),(2'd0)}}};
  localparam signed [4:0] p10 = {{(+(4'd7)),(^(3'd1))},((~|(4'd8))+(~^(-5'sd9)))};
  localparam signed [5:0] p11 = (((4'd0)|(2'sd1))>>((3'sd2)>>>(-4'sd6)));
  localparam [3:0] p12 = {((3'd0)==(3'sd3)),((2'd0)>>(3'd6))};
  localparam [4:0] p13 = {3{{4{(2'd3)}}}};
  localparam [5:0] p14 = (((5'd6)>(3'd0))?(-3'sd2):((-3'sd2)!=(3'd3)));
  localparam signed [3:0] p15 = (2'd3);
  localparam signed [4:0] p16 = ({((4'sd2)?(-4'sd6):(2'd0))}?((+(5'd3))&(|(5'sd2))):{(4'd4),(5'sd11),(-3'sd0)});
  localparam signed [5:0] p17 = {(~|(|{(~{(|(-4'sd4))}),(~((4'sd7)<<(-4'sd7))),(~&{(3'sd3),(4'sd7),(2'sd1)})}))};

  assign y0 = (+b4);
  assign y1 = (~|(3'd4));
  assign y2 = $signed((~^{(~{a2,b1,b4}),$signed(({b5,p5,b4})),((~|(~^(a0))))}));
  assign y3 = (|((!(|((p17<<p0)&(a3?p16:p2))))!=({4{a4}}?(+{p9}):(~^(p15?p1:p3)))));
  assign y4 = (2'd0);
  assign y5 = ((a3?a5:b1)?(-4'sd5):{{a3}});
  assign y6 = ({4{(a3?a5:a4)}}=={2{(~^{p11,b0})}});
  assign y7 = (((-3'sd0)>>(|p12))?(a4?a0:p0):((p17?p4:b0)>>>(4'd2 * p1)));
  assign y8 = (6'd2 * {4{a0}});
  assign y9 = ({4{{a5}}}>=(~(~^(5'd20))));
  assign y10 = (&(^a5));
  assign y11 = ({((b3<<p0)==(~p8))}>({p5,p9,p2}?{a3,p1}:(~&a0)));
  assign y12 = ((p14?p2:p8)?(p14?p6:p7):(2'd3));
  assign y13 = (~b5);
  assign y14 = ({2{b3}}?(p15):(p6));
  assign y15 = ({{b5,b3},(b2<=a4),(b4!==a2)}||{{b5},(a3===b5),(b1?b5:a4)});
  assign y16 = $signed(({1{b4}}-(b0==a4)));
  assign y17 = (~&(((~|(p1<<<p7))^((|p17)>>(p2&&p15)))>=((~^(~^(b5||p9)))|{(~&(!p1))})));
endmodule
