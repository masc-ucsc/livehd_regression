module expression_00292(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({((4'd1)===(4'd4))}?(!{4{(5'd23)}}):((3'd2)?(3'd6):(4'sd7)));
  localparam [4:0] p1 = (((-5'sd10)?(5'sd8):(3'sd3))?((3'd3)+(3'd6)):(~|((2'd0)?(5'd24):(2'd3))));
  localparam [5:0] p2 = {{(5'd2 * ((4'd12)&&(4'd15)))},((((3'd5)^(3'd6))-{(2'sd0),(-2'sd0),(2'd1)})!=(4'd2 * {(4'd8),(4'd3),(4'd13)}))};
  localparam signed [3:0] p3 = {2{{1{{4{(2'd2)}}}}}};
  localparam signed [4:0] p4 = {4{{(4'd9)}}};
  localparam signed [5:0] p5 = {2{{(^(~(((5'sd0)||(2'd0))&&(!(4'd15)))))}}};
  localparam [3:0] p6 = (({2{(3'd7)}}+(5'd21))?({(5'd28)}?((2'sd0)?(4'd6):(2'd1)):(~&(5'd9))):(2'd0));
  localparam [4:0] p7 = ({2{(5'd25)}}?(4'd15):(2'd2));
  localparam [5:0] p8 = {(((-3'sd2)|(-4'sd2))>>>{1{(&(3'd6))}}),({2{(4'd13)}}>>{3{(4'd13)}})};
  localparam signed [3:0] p9 = ((((3'd5)&&(5'd19))||{1{{(3'd4),(2'sd1)}}})<=({{(4'd7),(2'd1)}}||((3'sd2)<<<(2'd1))));
  localparam signed [4:0] p10 = ((((5'sd11)<<<(4'd3))?((3'sd1)?(2'sd1):(2'd3)):((5'd4)^~(5'sd1)))!==(((5'd26)>(-5'sd4))?(2'sd0):((3'd6)?(5'd30):(-4'sd2))));
  localparam signed [5:0] p11 = ((3'd1)?(&(-3'sd3)):((3'sd0)|(3'd7)));
  localparam [3:0] p12 = {{4{(-3'sd3)}},{1{{3{{2{(5'd18)}}}}}}};
  localparam [4:0] p13 = {3{(-2'sd0)}};
  localparam [5:0] p14 = (((|(3'sd2))<<((5'd13)===(4'd13)))||(((5'd6)^(-3'sd0))<(!(-5'sd9))));
  localparam signed [3:0] p15 = (~|(-3'sd0));
  localparam signed [4:0] p16 = (({(2'd1),(4'd0),(2'sd0)}-{(5'sd11),(2'd0),(3'sd1)})>({(3'sd0),(-2'sd0),(-2'sd0)}<=((3'sd1)==(2'd3))));
  localparam signed [5:0] p17 = (5'sd1);

  assign y0 = (~b4);
  assign y1 = {2{(+{4{p10}})}};
  assign y2 = (+{p10});
  assign y3 = {(|{(|(~a0))}),(^{p7,p3,b1}),{4{a4}}};
  assign y4 = {((-5'sd4)^{3{{3{p16}}}})};
  assign y5 = (~((a2?a1:p5)?(-4'sd1):(+(b1?p6:p3))));
  assign y6 = ((&((~^p12)?(p8?a4:a2):(-p4)))?({1{(-p3)}}&{4{a1}}):(~{3{(p2?p1:b0)}}));
  assign y7 = (({2{(a2===a5)}}|((b2?b2:b3)<<(b4>>a2)))<({3{(b3?p12:p12)}}&&{1{((p10<<b4)<=(p1>>>b0))}}));
  assign y8 = ((6'd2 * (+(3'd3)))?(-3'sd2):$unsigned(((!p1)?(p8?b3:p7):(~|p6))));
  assign y9 = (~&(4'd14));
  assign y10 = ((~(^(3'sd0)))|(-5'sd10));
  assign y11 = {4{(-4'sd3)}};
  assign y12 = {b3};
  assign y13 = (&(-4'sd2));
  assign y14 = (((2'd0)>=((p15<<p12)<<(-4'sd6)))<<<(~(~&(!((5'sd12)<(~|b0))))));
  assign y15 = ({3{{2{{2{b4}}}}}});
  assign y16 = (|((2'd1)<((~|(~^(+(a4*b5)))))));
  assign y17 = (!({(4'd2 * p14),(2'd3)}||(~^((p4+p13)>$unsigned(p2)))));
endmodule
