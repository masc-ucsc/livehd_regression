module expression_00727(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((4'sd6)?(5'd22):(-2'sd0)),((-2'sd0)&&(4'd3))};
  localparam [4:0] p1 = (({{(-3'sd2),(2'sd1),(5'd29)}}<=((5'd10)>(4'd8)))&(((-3'sd3)-(4'd6))^~((-5'sd9)<=(-5'sd14))));
  localparam [5:0] p2 = (({2{((4'sd7)&(3'd0))}}!==((-2'sd1)?(3'd2):(4'sd6)))&&({3{(-3'sd1)}}?{3{(2'd2)}}:((-5'sd3)||(2'd3))));
  localparam signed [3:0] p3 = ({(-2'sd1),(-2'sd0)}===(&(3'd3)));
  localparam signed [4:0] p4 = (+(~|(^(!(^(~(|(&(!(~(|(-5'sd12))))))))))));
  localparam signed [5:0] p5 = (-(+{2{(4'd2)}}));
  localparam [3:0] p6 = (+(2'sd1));
  localparam [4:0] p7 = (|(((-2'sd0)+(-3'sd1))!==(+((4'sd7)>>>(5'd17)))));
  localparam [5:0] p8 = ((5'd20)<<<(~^((~&(2'sd0))?((4'sd2)?(-4'sd0):(-4'sd5)):(~&(-4'sd1)))));
  localparam signed [3:0] p9 = (-(!(-(~&(&(+(&(^(!(~&(4'd11)))))))))));
  localparam signed [4:0] p10 = (((-3'sd1)?(3'd0):(4'd11))^((-4'sd3)?(2'd3):(-4'sd2)));
  localparam signed [5:0] p11 = (~|{((4'd4)<=(5'sd10)),((-5'sd8)^(2'd0)),{2{(3'd7)}}});
  localparam [3:0] p12 = ((5'd30)|(5'd2));
  localparam [4:0] p13 = {4{(2'd3)}};
  localparam [5:0] p14 = ({{(5'sd9),(5'd7),(-5'sd14)},({(3'sd1),(-5'sd5),(2'd0)}==((5'd27)<<(2'd1)))}<=((((-4'sd0)+(2'd0))<<((2'd3)<(5'd27)))+{(-5'sd12),(-3'sd1),(-5'sd12)}));
  localparam signed [3:0] p15 = (-4'sd4);
  localparam signed [4:0] p16 = (((4'sd2)?(2'd3):(3'sd0))+((3'd5)|(-2'sd0)));
  localparam signed [5:0] p17 = (2'd3);

  assign y0 = ({3{(a5||b2)}}>(&({1{(a3!==a1)}}^~{(a1<a2),{3{b1}}})));
  assign y1 = ({{2{b3}},{b2,b2}}?{2{{p11}}}:{1{(a2?p6:a3)}});
  assign y2 = ({2{(b1+a0)}}!==(5'd2 * (-a1)));
  assign y3 = {((b0?b0:p13)?{{4{b3}}}:{b0,b2,a0})};
  assign y4 = ((2'sd1)<<{{(b1==p12)},(p7&p13),(p5<<<a4)});
  assign y5 = (5'd18);
  assign y6 = {3{{2{(p9?b5:b2)}}}};
  assign y7 = ({p2,p8}>>(p2|p12));
  assign y8 = ($signed((&(-$unsigned((~^{(~&p14),(5'sd7),$unsigned(p6)})))))<<<$unsigned((-2'sd0)));
  assign y9 = {{2{({2{{a4}}}+{a0,b4,a0})}}};
  assign y10 = ((&(^(6'd2 * (4'd6))))-({3{a3}}>>>(|(5'd9))));
  assign y11 = {p9,p12,p15};
  assign y12 = (^((a2==a2)?(~^p8):(a5+a5)));
  assign y13 = (~&({a2,a4,b5}!==(b5?a3:a4)));
  assign y14 = (~&((((b1^~a2)<<(b2^a4))===((b0?a5:a4)!==(a4?b5:b1)))&(~^(!(~&(~&((p9<<p9)&(b4!==a3))))))));
  assign y15 = (-p15);
  assign y16 = {2{{2{(p6>>>p2)}}}};
  assign y17 = ({(a1?a0:b3),{a3,b3},(b5?b0:a4)}?((b5?b4:b5)?(&a4):(p7?a3:a1)):({b2}?(+a0):{a1,b2}));
endmodule
