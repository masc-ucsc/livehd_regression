module expression_00271(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'sd2)|(5'd16))-((-2'sd0)&(3'd5)))<=(((4'd15)==(-4'sd0))==((5'd10)&&(2'sd1))));
  localparam [4:0] p1 = (~&(~&(^(~&{(~{({(4'd12),(4'd0)}<<((-5'sd1)!==(-4'sd0))),{(5'd10),(5'sd12),(-5'sd6)}})}))));
  localparam [5:0] p2 = ({2{(-4'sd4)}}=={1{(-(-5'sd0))}});
  localparam signed [3:0] p3 = ((((-4'sd5)?(4'd0):(3'sd2))-((2'd3)?(5'd20):(-5'sd1)))!==(((-2'sd0)?(2'd1):(2'd0))==((-5'sd0)>>(-3'sd2))));
  localparam signed [4:0] p4 = ((-3'sd0)||(5'd23));
  localparam signed [5:0] p5 = ((5'd1)^~(5'sd5));
  localparam [3:0] p6 = (-4'sd3);
  localparam [4:0] p7 = {3{(-2'sd1)}};
  localparam [5:0] p8 = (+(|(-3'sd0)));
  localparam signed [3:0] p9 = ((~^((4'd13)?(4'd12):(-2'sd0)))===(~&((3'd6)?(4'd10):(3'd3))));
  localparam signed [4:0] p10 = ((((2'd1)^~(5'd4))|{4{(3'd5)}})>(((4'sd7)>(2'd3))^~((4'sd2)>=(2'd1))));
  localparam signed [5:0] p11 = (((6'd2 * (5'd10))<=((4'd10)?(2'd3):(5'd21)))?(!{(5'd2 * (2'd0)),((4'd1)^(-4'sd5))}):(((2'd2)+(-5'sd7))&(^(4'd9))));
  localparam [3:0] p12 = ((((5'sd8)?(5'd17):(2'd3))*((5'sd10)?(4'd8):(5'd20)))>(~^(((3'd5)?(-5'sd2):(2'd0))===((3'd1)?(3'sd2):(-5'sd8)))));
  localparam [4:0] p13 = (4'd11);
  localparam [5:0] p14 = ((-{((5'sd13)&&(-3'sd1)),(~(3'd5)),((-5'sd8)?(4'd4):(5'd17))})<(~|((~|(-4'sd0))&{(3'd6),(4'd4),(5'd19)})));
  localparam signed [3:0] p15 = (|{(~&(3'sd1)),(5'd2)});
  localparam signed [4:0] p16 = {(4'sd1),(2'sd1),(-5'sd2)};
  localparam signed [5:0] p17 = (~|(-4'sd5));

  assign y0 = (&(p5|a2));
  assign y1 = (-2'sd1);
  assign y2 = ((~|{4{(2'd1)}}));
  assign y3 = (^{1{{2{{2{a2}}}}}});
  assign y4 = $unsigned($unsigned($signed((-(~|(2'd3))))));
  assign y5 = (2'd2);
  assign y6 = ((~|((!(p3|p14))==((p11>p14)^~(p12<<<p7))))==({(p0?p3:p0),(p7<<b1)}==(~|(~^(5'sd12)))));
  assign y7 = (5'd28);
  assign y8 = ((-(~&(((|(~^b2))*(~(&p6)))))));
  assign y9 = $signed(({1{$signed(p9)}}==$signed((p1||p9))));
  assign y10 = {(2'd3)};
  assign y11 = (((p5-b0)?(b1<a3):(p11>>>a2))?({1{b3}}?(&b2):{p3}):{4{(~|a5)}});
  assign y12 = ((-(a2<<a0))>((&b3)&{a3,b5}));
  assign y13 = (|$unsigned((-(~|$unsigned((((p6?p15:p15)^~$signed(p4))?((p1<p8)|(p14?p17:p15)):((a3+a5)!==(b5||b5))))))));
  assign y14 = ((a5===b1)>>>(b0!==b0));
  assign y15 = (~|(5'd20));
  assign y16 = (-(|(((b4>>>a2)||(+(a1<b3)))&&{((a2===a0)&(|(!a5)))})));
  assign y17 = (~^(~&(!(-{1{{3{{3{{1{b5}}}}}}}}))));
endmodule
