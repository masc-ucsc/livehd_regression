module expression_00618(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{((4'd15)&&(-5'sd2)),((4'd7)>=(5'd17))},{(3'd5)}};
  localparam [4:0] p1 = {3{(+(-{4{(5'sd15)}}))}};
  localparam [5:0] p2 = (((4'd8)?(3'd4):(2'd2))^~((2'd1)?(2'd3):(-2'sd1)));
  localparam signed [3:0] p3 = (({(2'd2),(4'd14)}^~{(-4'sd5),(3'd7)})-(((4'd6)-(3'd7))^{(2'd2),(3'sd1)}));
  localparam signed [4:0] p4 = (+(-(-5'sd8)));
  localparam signed [5:0] p5 = (~|{3{({3{(4'd2)}}>>(^(-4'sd3)))}});
  localparam [3:0] p6 = (4'd10);
  localparam [4:0] p7 = ((|(2'd0))?((5'd19)?(4'sd4):(-2'sd0)):((4'd14)>>(5'd27)));
  localparam [5:0] p8 = (&(!(~^(!(~((|(&(5'd12)))>=(&(~(5'd29)))))))));
  localparam signed [3:0] p9 = ((-2'sd0)^~(3'd0));
  localparam signed [4:0] p10 = {{{(2'sd0),(2'd1),(2'sd1)},((2'sd1)?(3'd3):(2'd1)),((2'd2)^(3'd3))},(((2'sd1)?(-2'sd1):(-2'sd1))?((4'd0)>=(-5'sd3)):((5'd28)?(3'sd0):(5'd6)))};
  localparam signed [5:0] p11 = {3{(~&(4'd15))}};
  localparam [3:0] p12 = ({1{((2'sd0)<<(-5'sd13))}}!=={3{(-5'sd1)}});
  localparam [4:0] p13 = ((+((4'd7)?(3'd3):((2'd1)>=(2'd2))))&({4{(3'sd2)}}>>(|((5'sd9)?(2'd3):(3'sd3)))));
  localparam [5:0] p14 = {({4{(4'd14)}}+((4'd2)+(3'd5))),(((2'd0)!=(3'd2))>>((5'd11)&&(5'd3))),{{4{(2'd1)}},((-3'sd0)-(-4'sd0))}};
  localparam signed [3:0] p15 = ({(&(-5'sd2)),(|(2'd0))}&(+(5'd6)));
  localparam signed [4:0] p16 = (-5'sd2);
  localparam signed [5:0] p17 = (^(-((^((5'sd11)^~(4'd8)))*(~&((-2'sd0)-(5'd29))))));

  assign y0 = (~|((!(~&p16))%p11));
  assign y1 = (((4'd1)<={2{b1}})?{1{(5'sd13)}}:$unsigned(((2'd1)?$unsigned(a1):(p4<<b5))));
  assign y2 = $signed(((!(~&{p15,p10}))>=(~&$unsigned((p3)))));
  assign y3 = (((p0?p6:p1)+{1{(p16!=b2)}})<<(((~|p2)>>(p5^~b4))>(b0?b2:p17)));
  assign y4 = (~(a2>=b5));
  assign y5 = ((-({4{a1}}?(a2===b2):{a3,b2}))<<(~^((b2<<a1)===(a1>>a3))));
  assign y6 = (({3{b3}}?{3{a0}}:{a0,b4,a3})>((b4?b2:b0)+{(!{4{p2}})}));
  assign y7 = ((p10<<p12)+{4{p14}});
  assign y8 = ((a4?b5:a2)?(4'd11):(-2'sd1));
  assign y9 = (((p15?p13:p4)?(+p14):{1{p1}})?{2{(!{3{p0}})}}:(-4'sd1));
  assign y10 = {(5'd13),{(6'd2 * p7)}};
  assign y11 = {(~|{p13,a0}),(5'd5)};
  assign y12 = (^{2{(~|(~|(|(5'sd13))))}});
  assign y13 = (|(~&(&(((-(^(~&p6)))||{p11,b4,p5})||((p14?p12:a4)&&{(^p3),(+p17)})))));
  assign y14 = (&((p7?p16:p12)?(~&(p2?a0:p17)):(-(p13?p15:p2))));
  assign y15 = (6'd2 * (p8?b2:p0));
  assign y16 = ((2'd3)^(((~^b1)?(a1!==b2):(+b4))===((a1<=b1)?(~^b3):(b0?b4:a0))));
  assign y17 = {1{(^(((b2<=a1)<(~&p12))?((+p10)?(b1==b2):(b4>p6)):((p10-p2)<<<(+p10))))}};
endmodule
