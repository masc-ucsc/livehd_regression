module expression_00564(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd28);
  localparam [4:0] p1 = (-(((5'd19)>>>(3'd6))^(~((-4'sd1)*(3'd1)))));
  localparam [5:0] p2 = ((((2'd0)!==(3'd1))>>((2'sd0)+(5'sd4)))|(-4'sd0));
  localparam signed [3:0] p3 = {{(6'd2 * (5'd0)),((-4'sd7)>(3'sd0)),{(5'd22)}}};
  localparam signed [4:0] p4 = (((|(3'd3))|((2'd2)?(5'd15):(3'd3)))?(((2'd2)|(4'd13))?(2'd3):((2'd1)!=(-4'sd1))):(~^((3'd1)?(5'sd2):(4'sd4))));
  localparam signed [5:0] p5 = ((5'd25)!=(3'd0));
  localparam [3:0] p6 = (4'sd4);
  localparam [4:0] p7 = ((((5'd8)!==(-3'sd3))<(&(5'd5)))>=(|((~|(3'd7))<<(5'd9))));
  localparam [5:0] p8 = (2'd1);
  localparam signed [3:0] p9 = {1{({1{{((4'd4)>>(5'd4))}}}<<(-4'sd1))}};
  localparam signed [4:0] p10 = (({2{(3'd0)}}?{3{(5'sd13)}}:{3{(2'sd0)}})?{3{(5'd2 * (4'd8))}}:({1{(5'd20)}}-((5'd28)|(5'sd0))));
  localparam signed [5:0] p11 = ((3'sd2)?(4'd1):(3'sd0));
  localparam [3:0] p12 = (((5'd15)?(5'd21):(5'd18))?((-5'sd13)?(3'sd3):(2'd1)):((5'd17)?(5'd29):(3'd0)));
  localparam [4:0] p13 = ((&((|((2'd3)<=(4'd0)))==((4'd6)*(2'd2))))&((^(&(-4'sd7)))==((3'sd1)&(4'd8))));
  localparam [5:0] p14 = (-4'sd1);
  localparam signed [3:0] p15 = {(((3'd1)&&(4'd9))?((5'd17)!==(4'd13)):((-2'sd0)>>(-2'sd0)))};
  localparam signed [4:0] p16 = (5'sd6);
  localparam signed [5:0] p17 = {{(5'sd7),(4'd5)}};

  assign y0 = (((~|p0)<<<(!p10))?(^{(p0==p16),(+p0)}):((4'd2 * p8)?(-p13):{p3}));
  assign y1 = ((3'd2)>{2{(5'd29)}});
  assign y2 = {4{a1}};
  assign y3 = $signed((b4!=b2));
  assign y4 = {{p4,p14},(p17<<a4),(b0&&b3)};
  assign y5 = ($signed((~^(~(p2|p0)))));
  assign y6 = ((|(~^((a3^a2)&&(b1?p17:a4))))?((a0===a3)/b5):((&b4)?(a2?a4:b2):(a5>>>p9)));
  assign y7 = $unsigned((((b1||p0)==(p8?a1:p10))>>$signed($unsigned({p7}))));
  assign y8 = (((a4^~a5)?{a3,b0}:(+a1))^~((b5^a5)?(b4?p10:b1):(!b5)));
  assign y9 = $signed((+$signed(((^(~(4'd10)))))));
  assign y10 = ((p1==a4)/p8);
  assign y11 = (~{2{(p0^p11)}});
  assign y12 = ((p5<<<p10)?(2'd3):(2'd2));
  assign y13 = ({1{((b2?b3:a4)>>>({3{b4}}<<<(&a2)))}}==(((^a2)<<<(a0-b2))+((a0?a3:b2)==(a4^a5))));
  assign y14 = (2'sd0);
  assign y15 = ($unsigned(p8)>=(p0>>>a2));
  assign y16 = (((a2===a2)<<<(p8?p5:p3))^((2'd2)?(3'd7):(p7?a4:p13)));
  assign y17 = (5'd2 * (+{2{a1}}));
endmodule
