module expression_00751(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd0)};
  localparam [4:0] p1 = {(-2'sd1),(((-4'sd1)?(3'sd3):(-2'sd1))?(^(-5'sd10)):(^(2'd0))),(^(4'd8))};
  localparam [5:0] p2 = ((3'sd3)<<((3'sd0)^(3'd7)));
  localparam signed [3:0] p3 = ((4'd13)+{2{{1{(-2'sd1)}}}});
  localparam signed [4:0] p4 = (((3'd3)%(2'sd1))*(5'd2 * (5'd19)));
  localparam signed [5:0] p5 = ((((5'd10)-(5'd17))||((4'd12)&&(5'd5)))+(((2'd1)>>(-3'sd1))<<((4'd12)^(4'd0))));
  localparam [3:0] p6 = ((&(!(-4'sd5)))||((-2'sd1)&(2'd0)));
  localparam [4:0] p7 = {{4{{3{(4'd13)}}}}};
  localparam [5:0] p8 = ((((5'sd11)|(3'sd2))!==(5'd2 * (2'd1)))!==(~&(~(+(~|((2'sd1)||(3'sd0)))))));
  localparam signed [3:0] p9 = (!{{(-4'sd3)},(~(5'sd10))});
  localparam signed [4:0] p10 = (^(~&{{(5'sd8),(4'd0),(-5'sd13)}}));
  localparam signed [5:0] p11 = (&(5'd3));
  localparam [3:0] p12 = ((((3'sd3)>=(3'd0))&((-2'sd0)===(2'd1)))<={3{{(4'd2),(5'd15)}}});
  localparam [4:0] p13 = (~^(({2{(3'd1)}}?(4'd2 * (3'd0)):{1{(3'd0)}})>>{3{(!(3'd6))}}));
  localparam [5:0] p14 = (4'd2 * ((3'd6)||(3'd0)));
  localparam signed [3:0] p15 = (3'd0);
  localparam signed [4:0] p16 = (&((4'sd6)==(-2'sd1)));
  localparam signed [5:0] p17 = {{{(2'd0),(2'd0)},{(-3'sd2)}},{(!(-4'sd4)),(|(3'd6))}};

  assign y0 = {((^(&(p2>=b0)))<<{(|{1{(b3?b5:a3)}})}),({3{p4}}?(a1!==b4):(p13?a4:p8))};
  assign y1 = $signed((^(-3'sd2)));
  assign y2 = {3{{2{{2{p16}}}}}};
  assign y3 = (({4{p11}}<=((b5>>a0))));
  assign y4 = (((a0?p9:p0)?(b2?p10:b2):(+p12))-(~|(~^{4{b2}})));
  assign y5 = (~|((-(3'sd1))^~(-((|{1{b5}})!=(+(2'd2))))));
  assign y6 = ((b0!==a4)+{1{b2}});
  assign y7 = {2{p12}};
  assign y8 = {1{((b0^p3)==(&p15))}};
  assign y9 = ((($signed(p11)|(p7?p6:p2))<((p0+p15)-(b1||p0))));
  assign y10 = ((2'd2)?(p13>p15):(-2'sd0));
  assign y11 = ($signed($signed(((&(b5||a4))&&(a5<b0))))===(((b4)&(a0===a4))>=((b2)&(b0==a5))));
  assign y12 = ({(5'sd4),(3'd7)}=={(5'd2)});
  assign y13 = (|p4);
  assign y14 = (({4{b2}}?{a3,b3,a0}:(a2?a5:p16))<<{(b1>p5),(p2?p3:p1),{b5,p12,p14}});
  assign y15 = (((p0|a1)<(p14==p2))?((2'sd1)<<{1{(p17?p13:b3)}}):($unsigned((a2?a2:a1))>>>(a1===b3)));
  assign y16 = ({4{(p17|b5)}}+{{b0,a3,b3},{4{b5}},(a1>=a3)});
  assign y17 = (2'd3);
endmodule
