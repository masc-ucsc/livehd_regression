module expression_00581(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'sd0)!==(-2'sd0));
  localparam [4:0] p1 = (5'd4);
  localparam [5:0] p2 = ({1{(-(4'd13))}}<=(^{1{(5'd24)}}));
  localparam signed [3:0] p3 = (3'd4);
  localparam signed [4:0] p4 = (((2'd1)?(4'd5):(4'sd7))?((-5'sd12)?(2'd2):(5'd25)):((3'd3)?(2'd3):(2'd2)));
  localparam signed [5:0] p5 = (|(&(~^(~(~|(^(5'sd1)))))));
  localparam [3:0] p6 = {3{(&(-4'sd3))}};
  localparam [4:0] p7 = {1{(~^(((4'd14)?(5'd23):(2'd2))?((5'sd10)?(5'd15):(2'd3)):((2'd0)?(2'd0):(2'd3))))}};
  localparam [5:0] p8 = ((-2'sd0)?{(2'sd1),(5'sd6),(-5'sd1)}:(+(3'sd2)));
  localparam signed [3:0] p9 = (~|{((5'd10)+(2'd2)),(^{(3'd3)}),{(2'sd0),(5'sd4)}});
  localparam signed [4:0] p10 = (({1{(3'sd2)}}+((4'sd6)!==(2'sd0)))==(((-5'sd12)?(-3'sd2):(3'd7))||{3{(2'd2)}}));
  localparam signed [5:0] p11 = (((~^((4'd7)>=(4'd5)))>>>((3'd7)^(3'd5)))-({(-5'sd7),(3'd6)}+{(2'sd1),(4'd3),(4'sd4)}));
  localparam [3:0] p12 = (~((4'd2)|((2'd1)>>>(-3'sd0))));
  localparam [4:0] p13 = (-(4'sd4));
  localparam [5:0] p14 = (((-3'sd3)?(4'd1):(2'd0))?((4'd15)^~(-4'sd5)):((-2'sd0)|(2'd1)));
  localparam signed [3:0] p15 = ({3{(2'd2)}}^~{2{(2'd2)}});
  localparam signed [4:0] p16 = (((-3'sd1)||(5'd0))=={4{(5'd16)}});
  localparam signed [5:0] p17 = {1{(((3'd7)<(-4'sd6))===(-5'sd2))}};

  assign y0 = (((!(a4?p5:b5))?{a1,a2}:(~^(a3^a0)))<(&(-((6'd2 * b2)?(p9&a1):(b0+b0)))));
  assign y1 = ({a4,a5,p5}>>(&p10));
  assign y2 = $signed($signed((2'sd1)));
  assign y3 = {{(p7==b0)},{{p10,p11,p10},(-p1)},(^(p11==p12))};
  assign y4 = (((p3?a4:p0)==(-(p2^p15)))==$unsigned((~|((p9?p17:a1)))));
  assign y5 = {{(({p7,p14}||(a5>>>b5))+((p10|b1)-{p17,b3})),({{b2,p3},(p1>>a5)}^({p4,p16}<<<{b0,p14}))}};
  assign y6 = (^(&(-2'sd0)));
  assign y7 = (4'sd7);
  assign y8 = (((|b4)));
  assign y9 = (+((($unsigned(a5))>>>(a0/b3))-$signed(($signed((b2||b3))%a4))));
  assign y10 = (~|$signed((3'sd1)));
  assign y11 = (((b1||b0)?(b1?a1:p3):{3{a1}})^({2{(a4|b0)}}>>((b2-b3)?(a4?b0:a0):(a2>>a1))));
  assign y12 = (4'd2 * (b2===a2));
  assign y13 = {({(5'd5),(3'd6),(p2==p6)}<{3{{p12,p0}}})};
  assign y14 = ((p7?a3:b0)?(b0?b5:b2):{(b3?b2:a2),{a1}});
  assign y15 = {1{(~|(-(~&{2{(~(^a1))}})))}};
  assign y16 = $unsigned((~&$unsigned((($signed((4'd2 * a2))!==(&(&a4)))))));
  assign y17 = (4'sd6);
endmodule
