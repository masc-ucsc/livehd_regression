module expression_00463(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^{(3'sd0)});
  localparam [4:0] p1 = (^((!(2'sd1))>=(+(2'd2))));
  localparam [5:0] p2 = (-3'sd2);
  localparam signed [3:0] p3 = (-(((4'd1)+(-4'sd4))/(5'd28)));
  localparam signed [4:0] p4 = ((((4'sd3)&&(2'd1))^~((4'd8)==(2'd0)))<=((&((3'sd1)>=(4'd5)))<(4'd2 * (5'd15))));
  localparam signed [5:0] p5 = ({(4'd3),(5'd14),(2'sd0)}?({(4'sd4),(4'sd4)}>>>((2'd3)?(-3'sd2):(2'sd1))):((3'd3)?(-2'sd1):(-3'sd2)));
  localparam [3:0] p6 = (((-5'sd4)>>>(-2'sd1))>>(-3'sd3));
  localparam [4:0] p7 = (^(-(((-3'sd2)|(-5'sd5))<=(-3'sd0))));
  localparam [5:0] p8 = (-((&(3'sd3))&&(!(2'd1))));
  localparam signed [3:0] p9 = {((2'd0)?(4'd3):(5'd30)),{((4'd6)?(4'd2):(4'd3))},((2'sd0)?(5'sd12):(2'd2))};
  localparam signed [4:0] p10 = ((((2'sd0)&(-2'sd0))<=((2'sd1)==(-4'sd1)))<<<(((2'sd0)==(-4'sd0))!==((3'd6)-(2'd2))));
  localparam signed [5:0] p11 = (((3'd1)<((3'sd1)<<(2'd2)))!==(|(((4'd15)?(3'd1):(3'd7))?((2'd3)*(5'd27)):((5'sd11)>=(5'd27)))));
  localparam [3:0] p12 = ((-4'sd6)&(5'sd7));
  localparam [4:0] p13 = ((-2'sd0)?{1{(5'd20)}}:(2'd1));
  localparam [5:0] p14 = ((3'sd0)<<<(4'sd0));
  localparam signed [3:0] p15 = ((5'sd13)!==(-3'sd0));
  localparam signed [4:0] p16 = ({4{(3'd6)}}===(2'd0));
  localparam signed [5:0] p17 = (3'd7);

  assign y0 = ((p4>>>a0)?(b5?p15:b0):(b4?a3:a2));
  assign y1 = (~&((3'd5)!=={{b4,b5,a0}}));
  assign y2 = (b1^a2);
  assign y3 = {(~|(-2'sd0))};
  assign y4 = ((-3'sd1)%a2);
  assign y5 = (|((p6+p8)));
  assign y6 = {2{{2{p1}}}};
  assign y7 = {(2'd3),(-2'sd0)};
  assign y8 = ((p15?p12:b2)||((p4>p6)));
  assign y9 = {($unsigned((2'sd0))),$unsigned($unsigned((4'd8))),{($signed({a5,b0,b3}))}};
  assign y10 = {$signed((({p15}?(b1<<<a0):{b3}))),((b5<<<a0)?(~&(a4)):$unsigned($signed(a2)))};
  assign y11 = (3'sd3);
  assign y12 = {a2,a0};
  assign y13 = {3{$signed(p3)}};
  assign y14 = $unsigned((-(^{$unsigned(($signed(((&((-{{a2,a3,a0},(^{b2}),$signed($unsigned(a2))})))))))})));
  assign y15 = {2{(5'd2 * (b1>p13))}};
  assign y16 = (~&(3'd2));
  assign y17 = (5'd27);
endmodule
