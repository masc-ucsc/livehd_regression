module expression_00298(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'd8);
  localparam [4:0] p1 = (^(|(-5'sd2)));
  localparam [5:0] p2 = (5'sd5);
  localparam signed [3:0] p3 = (((!(3'sd0))>=((5'd20)?(4'sd6):(2'd1)))&&((~&(2'd3))?(-(-5'sd4)):((4'd0)!=(5'd21))));
  localparam signed [4:0] p4 = ((&(^((4'd4)^(3'sd3))))?(((-3'sd2)?(5'd31):(2'd2))&((5'd7)?(5'sd6):(-5'sd7))):(&(~&((3'd7)?(4'd8):(-2'sd1)))));
  localparam signed [5:0] p5 = (!{((-2'sd1)>(((4'd13)>>>(4'd10))&&((2'd0)<(5'd19))))});
  localparam [3:0] p6 = (~|{3{(2'd1)}});
  localparam [4:0] p7 = ((5'sd15)*(-5'sd15));
  localparam [5:0] p8 = {1{{3{(((2'sd1)<<<(2'sd1))!==((3'sd1)>>(5'd5)))}}}};
  localparam signed [3:0] p9 = ({{1{(-3'sd1)}},{(5'd12),(4'd11)},((-5'sd1)<<(5'd24))}<<<{3{(5'sd2)}});
  localparam signed [4:0] p10 = (~^(-3'sd0));
  localparam signed [5:0] p11 = (((-3'sd2)>(3'd0))+{(3'sd3)});
  localparam [3:0] p12 = {(((2'sd1)!=(-2'sd0))>>{(-5'sd0)}),((-5'sd15)+((5'd21)+(3'sd1))),(6'd2 * {{(4'd12),(5'd27),(4'd4)}})};
  localparam [4:0] p13 = ((5'sd0)?(4'd0):(4'sd0));
  localparam [5:0] p14 = (3'd5);
  localparam signed [3:0] p15 = (~&(-3'sd2));
  localparam signed [4:0] p16 = (((5'sd1)<<<(2'd0))?((-4'sd4)?(-3'sd3):(4'sd4)):((3'sd3)===(4'd7)));
  localparam signed [5:0] p17 = {{4{(&{(|(-4'sd0))})}}};

  assign y0 = (((a2^~b5)&&((b5<=b1)))||{{p13,a5,a0},(a0?b0:b2)});
  assign y1 = (~^((|(-(+p5)))));
  assign y2 = (2'd3);
  assign y3 = $signed($unsigned((-(^(2'd3)))));
  assign y4 = (~^(^(3'sd0)));
  assign y5 = (~(|$unsigned((~|(4'd5)))));
  assign y6 = (|{(5'sd12)});
  assign y7 = (!$unsigned(((~^($unsigned((p12&&b4))<(~(p11<<p10)))))));
  assign y8 = (2'd3);
  assign y9 = (((-3'sd3)/p17)!=(4'd10));
  assign y10 = {2{((p13)<<<(b3!==b1))}};
  assign y11 = (-4'sd0);
  assign y12 = (-4'sd5);
  assign y13 = (^{(|(&((p14?p6:p14)&(p8^p5))))});
  assign y14 = ({b0,a3}?(&(b4?b1:p11)):{a0,p9,p17});
  assign y15 = $signed({$unsigned((((b3<a3)+{b3,b4})|$signed(((b2|b4)!=(a3?b1:b5)))))});
  assign y16 = (!$unsigned((~^(~|$unsigned(((p15>=p13)!=(~^b0)))))));
  assign y17 = (-(!{2{(|{4{a3}})}}));
endmodule
