module expression_00941(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd2)<<(2'sd1));
  localparam [4:0] p1 = {{3{(!(-2'sd0))}},{(~|(4'sd7))},{2{(+(2'd3))}}};
  localparam [5:0] p2 = (-(5'd2 * ((3'd4)==(3'd0))));
  localparam signed [3:0] p3 = ((-3'sd1)||((^(4'd6))+((2'd2)>>(-4'sd1))));
  localparam signed [4:0] p4 = (4'd5);
  localparam signed [5:0] p5 = (-3'sd0);
  localparam [3:0] p6 = (&(-3'sd3));
  localparam [4:0] p7 = (-(((4'd3)?(5'd25):(3'd7))&((-2'sd1)>>>(3'd3))));
  localparam [5:0] p8 = {2{((4'd2 * (3'd0))?(5'sd13):{3{(2'sd1)}})}};
  localparam signed [3:0] p9 = (((4'd2)/(-2'sd1))>=(&(+(-3'sd0))));
  localparam signed [4:0] p10 = (+(((^(3'd7))<<<((3'sd1)>(5'd0)))||(+{(-4'sd2),(4'd10)})));
  localparam signed [5:0] p11 = ((((3'sd3)?(4'd14):(2'd3))?((5'd11)?(4'd12):(3'd6)):((4'd7)?(5'd25):(4'd11)))?(((4'sd0)?(3'd4):(4'd10))?((4'sd4)?(3'd6):(-2'sd1)):((-2'sd0)?(5'd18):(-4'sd6))):(((5'd0)?(3'd6):(-5'sd0))?((-4'sd4)?(-5'sd14):(5'd31)):((2'sd0)?(-4'sd2):(-3'sd3))));
  localparam [3:0] p12 = ((5'sd11)?{((-4'sd6)?(3'd4):(5'd9))}:(((3'sd1)<<<(4'd8))?(&(5'd1)):((-4'sd7)===(4'sd1))));
  localparam [4:0] p13 = ((^(~(+(!(5'sd13)))))?(^(-(&((5'd29)?(2'sd0):(2'd3))))):(~|(~&((5'd17)?(4'd14):(5'd10)))));
  localparam [5:0] p14 = ((~|(~|(2'sd1)))/(-3'sd2));
  localparam signed [3:0] p15 = (~|(-(((2'sd1)?(4'sd2):(4'sd3))^{(3'd1),(2'sd1),(4'sd5)})));
  localparam signed [4:0] p16 = {(3'd4),(-2'sd1)};
  localparam signed [5:0] p17 = (6'd2 * (5'd5));

  assign y0 = (!{3{(3'd4)}});
  assign y1 = (2'sd1);
  assign y2 = (~&(|(~&{(b3?p5:p1),(+(b5!==a2)),(p16|b4)})));
  assign y3 = ((p14&&p9)?(p3/p1):(p4?b5:p12));
  assign y4 = (|(a0===a5));
  assign y5 = ((a3?a4:a5)^~(a2+b5));
  assign y6 = ((b1?b0:b5)>>>{a3,p0,p0});
  assign y7 = (p5|p11);
  assign y8 = (^((b3-p13)+(a1?p16:p17)));
  assign y9 = ((p1<p11)?{1{(p4<=p10)}}:(p7<p4));
  assign y10 = {((($signed((a0?b5:a1))?(b4^~a1):{a4,b0,a1})>=({$signed(a4)}?($unsigned(b0)):$unsigned((p13?a1:p6)))))};
  assign y11 = (-(+(~&(~^(~|(!(!(~(~&(|(~^p7)))))))))));
  assign y12 = $unsigned($unsigned({4{$unsigned(a1)}}));
  assign y13 = (((!(a0>=a3))>>>((a1?a5:b4)&&(b5^~b5)))!==(~^(((+b0))==(b2?a2:a3))));
  assign y14 = {1{((b0?a2:a0)>>>(b2^~b4))}};
  assign y15 = (((b0?a5:p0)?$signed(b3):(!b3))?(&(p1?p9:a0)):(-($unsigned($signed(a0)))));
  assign y16 = {2{(3'd7)}};
  assign y17 = (p0-p5);
endmodule
