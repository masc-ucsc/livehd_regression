module expression_00886(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd4)?(-4'sd4):(5'd18))?((4'sd3)?(5'd9):(3'd3)):((-2'sd0)?(-3'sd1):(-5'sd12)));
  localparam [4:0] p1 = ((((2'sd1)<(3'sd2))>=(5'd2 * (2'd0)))>=({3{(3'sd1)}}+((-3'sd3)+(5'd20))));
  localparam [5:0] p2 = {{((-2'sd1)?(5'd31):(3'd6))},({(5'd21),(-4'sd5),(-2'sd0)}?(2'd2):((4'sd4)?(4'd5):(3'sd3))),(-2'sd0)};
  localparam signed [3:0] p3 = {3{{4{(3'sd3)}}}};
  localparam signed [4:0] p4 = {1{((+(|{1{({3{(2'sd0)}}^~(~^(2'd2)))}}))&&(|{4{{2{(5'd17)}}}}))}};
  localparam signed [5:0] p5 = (|(!(((2'd1)<<<{(-4'sd0),(-3'sd3),(3'sd2)})>>>(5'd2 * (+(2'd0))))));
  localparam [3:0] p6 = (5'sd11);
  localparam [4:0] p7 = (~|(^((&(5'd13))>=(^(2'd3)))));
  localparam [5:0] p8 = (5'd28);
  localparam signed [3:0] p9 = ((^((-5'sd8)>>>(2'sd0)))-((-2'sd0)&(5'sd10)));
  localparam signed [4:0] p10 = (-((4'd7)?(-2'sd1):(-3'sd1)));
  localparam signed [5:0] p11 = {3{((2'sd1)===(4'd4))}};
  localparam [3:0] p12 = {({(3'd1),(-2'sd0),(2'sd1)}-((3'sd1)?(4'sd3):(2'd1))),((-5'sd1)?(2'sd1):(5'sd8)),((-4'sd0)>(5'd14))};
  localparam [4:0] p13 = (-({1{(!((-2'sd0)>>>(2'd1)))}}<<(!{(-5'sd5),(-5'sd1),(3'd0)})));
  localparam [5:0] p14 = ((3'd6)?(2'd2):(4'd0));
  localparam signed [3:0] p15 = (&(^(|(~(5'd2)))));
  localparam signed [4:0] p16 = ((3'd3)?(-3'sd0):(3'd7));
  localparam signed [5:0] p17 = ((-2'sd0)?(3'sd2):(-3'sd0));

  assign y0 = {(^(-b1)),(p6?p7:b1)};
  assign y1 = {(-((p9>>>a0)<=(5'd20))),(4'd12)};
  assign y2 = (-(~&(!(p5|p4))));
  assign y3 = (~^((^(a4==b1))|(p16?a0:b2)));
  assign y4 = {{{p15,a5,p4},{(b1>>a3)},{p1,p14,p7}},{((p16<<a5)+(a5===a4)),({p1,p9}>{a5,p2})}};
  assign y5 = $signed($signed((a1|a0)));
  assign y6 = (+(((~|(~|(b0))))!==((~b5)|$unsigned(b2))));
  assign y7 = (5'd2 * (p0?p6:p6));
  assign y8 = {b3,a4,a1};
  assign y9 = (2'd0);
  assign y10 = ((-(~((p0?p3:p3)?(5'd1):(4'd9))))?(!((-2'sd1)?(&b3):(2'sd1))):((-3'sd3)?(~p17):(+a0)));
  assign y11 = {4{$signed($signed({1{p8}}))}};
  assign y12 = (~&(4'sd7));
  assign y13 = $signed((&{(!(b2?p12:b1)),(+$signed((3'sd3))),(+(4'sd6))}));
  assign y14 = ({2{(2'd1)}}?(-4'sd4):(^(^(b2?b3:b3))));
  assign y15 = (~&(&((5'd24)<=(+{(p17==p13),(~&p2),(+p2)}))));
  assign y16 = (($signed($unsigned((a3|b2)))>>((^b2)&(|b2)))!==(((b3&b5)+(a3||a2))>>>($signed(b0)!==(&a1))));
  assign y17 = (($signed((&(&(!((~p8))))))));
endmodule
