module expression_00579(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(((-5'sd13)===(-3'sd0))*((5'sd0)>=(4'd10))));
  localparam [4:0] p1 = (~&(-4'sd4));
  localparam [5:0] p2 = {(((-3'sd0)&&(3'sd3))?(^(-3'sd2)):(^(4'd1)))};
  localparam signed [3:0] p3 = {2{((5'd23)==(4'd11))}};
  localparam signed [4:0] p4 = {({(4'd12),(5'sd11)}!==(~(5'sd6))),(3'd6),{(4'd10),(3'd6),(3'd4)}};
  localparam signed [5:0] p5 = (((5'd4)?(4'd10):(2'sd1))^~{(2'd2),(5'sd14),(-4'sd3)});
  localparam [3:0] p6 = (({(!(3'd3))}|{(5'd31),(-2'sd1)})&&(-{(4'd2 * (-(-(3'd1))))}));
  localparam [4:0] p7 = ((((5'd1)<<<(-2'sd1))?((2'sd0)?(2'd2):(2'd2)):((-5'sd15)?(-2'sd1):(-5'sd6)))|((~&((5'sd3)/(3'd0)))&&(~&(!(2'd1)))));
  localparam [5:0] p8 = {(4'd12),(4'sd0)};
  localparam signed [3:0] p9 = (|({(((-3'sd3)&(4'd3))&(|((5'sd4)>>>(3'd6))))}<(+{1{(~|((^(3'sd3))+{(3'd1)}))}})));
  localparam signed [4:0] p10 = ({2{(5'd20)}}===(|(3'd5)));
  localparam signed [5:0] p11 = (((5'd20)!=(4'd7))*(|(2'd3)));
  localparam [3:0] p12 = (&((((-3'sd3)||(-5'sd13))>>>((2'd1)||(3'd7)))>>{(((-4'sd6)-(4'sd3))<<((5'd25)^(2'd0)))}));
  localparam [4:0] p13 = ((2'd3)!==(4'sd5));
  localparam [5:0] p14 = (((-2'sd0)<<<{4{(5'd8)}})&&((-4'sd0)<=((5'd4)===(4'd7))));
  localparam signed [3:0] p15 = (3'd6);
  localparam signed [4:0] p16 = (3'd5);
  localparam signed [5:0] p17 = {(~|((((-3'sd3)?(4'sd1):(2'd0))+((-4'sd7)?(-3'sd0):(-3'sd2)))>=(((4'd11)^(-3'sd0))?((-4'sd5)?(5'd3):(3'sd1)):((4'd8)!==(3'd2)))))};

  assign y0 = (~(a3?p15:p7));
  assign y1 = ((6'd2 * {p6,p0})&&{(p13^a1),{(p11<<p3)}});
  assign y2 = (~&(((a2?p5:b5)<=(~|b3))>=((b0?a3:p13)?(b5?b0:p3):(a0?a1:b2))));
  assign y3 = ((b1?p9:p5)<<{p2});
  assign y4 = (~&{($unsigned((!b5))),{{p5,b4}}});
  assign y5 = ((a0?a5:b2)===$unsigned((a2?a5:a5)));
  assign y6 = ((p10?p16:p4)?(p15?p15:p11):(|p16));
  assign y7 = (((p11<<<a1)>(b3&&a0))<<(~^((3'd3)==(-{b5,b2}))));
  assign y8 = (3'sd3);
  assign y9 = (!((~{1{({4{p4}}!={1{(a0||a0)}})}})^~{1{((~^{1{{4{p14}}}})||(+{1{{4{a1}}}}))}}));
  assign y10 = ((($signed(p4)+(4'sd7))&&{p12,p4,p17})==((4'sd5)==((a1<<a4)!==(b5==a3))));
  assign y11 = (p11?p15:a4);
  assign y12 = ({3{(-(|a4))}}-(|{2{((a4&a4)^(b3<<b4))}}));
  assign y13 = {b2,p10};
  assign y14 = ((~&{2{(4'sd7)}})&&(~(~|(~|(~|(~|{1{{3{p0}}}}))))));
  assign y15 = (5'd11);
  assign y16 = (~&({((~(~&b4))||(b0>>a4))}==({(b5<<<b0),{b2,a5,a4}}==(^{a2,a4}))));
  assign y17 = (^(+((2'd1)?((b2?p11:p17)^~$signed((5'd2 * a0))):((a4!==a1)<<<(p5>=a4)))));
endmodule
