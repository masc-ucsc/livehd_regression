module expression_00343(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-{3{((5'd20)>>>(2'sd0))}});
  localparam [4:0] p1 = ({2{(3'd3)}}>>>{4{(2'd0)}});
  localparam [5:0] p2 = ((-{3{{4{(5'd10)}}}})<<(((2'sd1)<<(-3'sd0))>>(^(~&(2'd3)))));
  localparam signed [3:0] p3 = (((-5'sd7)-((4'd10)>>(4'sd7)))>(~|(-5'sd1)));
  localparam signed [4:0] p4 = (5'd6);
  localparam signed [5:0] p5 = (-(^(~((2'sd1)?(2'd1):(3'd2)))));
  localparam [3:0] p6 = (((-2'sd0)>>>(3'd7))?(2'd0):(&(~&(2'd2))));
  localparam [4:0] p7 = {2{{4{(-2'sd1)}}}};
  localparam [5:0] p8 = ((((3'd6)&(3'd3))?(2'sd1):((2'd1)&&(5'sd15)))<(((2'd2)?(4'd11):(5'd31))&&((-2'sd1)!=(-3'sd2))));
  localparam signed [3:0] p9 = (~&{{{(2'd0),(-5'sd1),(4'd6)},{(3'd6),(2'd3),(4'sd4)},{(-4'sd1),(4'd6)}},({(5'd11),(3'd7),(2'd0)}!==((-4'sd0)^(2'd1))),{((-3'sd1)&&(2'd3)),{(3'd3),(3'd7)}}});
  localparam signed [4:0] p10 = ({{3{(2'd3)}},{(5'sd11),(-5'sd13)},(6'd2 * (2'd2))}&(~&{((4'sd1)<<<(5'd31)),((5'd24)&&(2'd1)),{3{(2'd0)}}}));
  localparam signed [5:0] p11 = (+(((-4'sd6)?(-5'sd7):(5'd9))^~(((2'sd0)!=(-3'sd1))^~{(3'd6)})));
  localparam [3:0] p12 = ((&{1{((4'sd6)+(-5'sd13))}})===(((2'd3)|(3'd2))!=(|(4'd9))));
  localparam [4:0] p13 = (3'd7);
  localparam [5:0] p14 = ((-3'sd0)?(-3'sd0):(5'sd8));
  localparam signed [3:0] p15 = (6'd2 * ((4'd4)^(4'd2)));
  localparam signed [4:0] p16 = (~&(6'd2 * (3'd2)));
  localparam signed [5:0] p17 = (((2'sd1)<<(-5'sd5))<=(-((-5'sd1)^(-2'sd0))));

  assign y0 = ((-$unsigned((~|$unsigned(a1))))>>>(~{1{(+(4'd2 * p2))}}));
  assign y1 = $unsigned(((((b3<a4)?(b5%a4):(^a3)))||((a0?b3:a4)?(b3?a0:b2):$unsigned(b3))));
  assign y2 = ((p15+p16)+{b3,p17,p6});
  assign y3 = ({$signed(p11),(6'd2 * p14)}&((p12&p13)+$unsigned(p0)));
  assign y4 = (|(((($unsigned(b1)?(p1>>>b5):$unsigned(a5))>((^a3)^(^b1))))));
  assign y5 = ($unsigned($unsigned($signed($unsigned(p5))))<<<((a3<b5)<<(2'd3)));
  assign y6 = (2'd1);
  assign y7 = $unsigned((((b2*b5))/a1));
  assign y8 = (((+p5)<(b1?p2:a2))^~(|(^(p3&b1))));
  assign y9 = {4{(!(-2'sd0))}};
  assign y10 = ((p13&p3)&(2'd3));
  assign y11 = ((a0?b3:p7)<(p8+p5));
  assign y12 = (b1<a2);
  assign y13 = ((((|p8)>>(p16&&a1))<<<$unsigned(((|a0))))>=(!((!(a3*p15))>>(-(a3-b0)))));
  assign y14 = {{p8,p5,p5},(p7^a4),(a3===a2)};
  assign y15 = (!((5'sd13)?((b0?p8:p6)|(a5?p15:p17)):((p4<p4)<(2'd0))));
  assign y16 = ((&((&(b3^~b2))>>>(&(a1%p5))))&((~(p8?a1:a2))<<<((~&p16)?(!p5):(|a0))));
  assign y17 = (((+(p12%p5))+(b5!==b5))<<(~|(|(a4?b3:a3))));
endmodule
