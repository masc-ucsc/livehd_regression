module expression_00412(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~((3'd0)<(3'd7)))<=((~^(-2'sd1))<((2'd0)<<(-4'sd4))))&((+((3'd6)-(-2'sd1)))&&((~(4'd9))-(|(4'd8)))));
  localparam [4:0] p1 = {(~(5'd25)),{(4'sd2),(4'sd2),(5'd27)}};
  localparam [5:0] p2 = (((5'sd13)?(3'd7):(3'd4))?((4'sd0)?(-3'sd3):(3'd5)):((-4'sd2)?(4'd0):(5'd9)));
  localparam signed [3:0] p3 = {3{{1{{4{(3'sd2)}}}}}};
  localparam signed [4:0] p4 = ((!(|(5'd2)))&&(4'sd1));
  localparam signed [5:0] p5 = {(3'd4)};
  localparam [3:0] p6 = (!(&{(-2'sd0),{(-4'sd0),(3'sd0),(2'd1)},{(4'd15),(4'd4),(-3'sd0)}}));
  localparam [4:0] p7 = (^{4{(2'd1)}});
  localparam [5:0] p8 = (5'd13);
  localparam signed [3:0] p9 = (-((-4'sd6)===(4'sd0)));
  localparam signed [4:0] p10 = {(5'd15),{(4'd15),(-5'sd4)},(4'd11)};
  localparam signed [5:0] p11 = ({1{((3'd4)?(4'd5):(-3'sd1))}}?(((5'd27)!==(2'sd0))<<((4'd11)?(2'd1):(2'sd1))):({1{(4'd13)}}|((2'sd0)+(5'd3))));
  localparam [3:0] p12 = {(+((5'd23)?(-2'sd0):(2'd1)))};
  localparam [4:0] p13 = {(~(2'd0))};
  localparam [5:0] p14 = {2{((3'd4)<<(2'd2))}};
  localparam signed [3:0] p15 = ((~(~^(((5'sd11)^~(4'd14))?((3'd2)|(5'd23)):{(4'd8),(4'd3)})))^~(3'd0));
  localparam signed [4:0] p16 = (~|((^{4{(4'd2)}})&&((-4'sd3)^~(-3'sd0))));
  localparam signed [5:0] p17 = ((+(4'sd0))<((4'd7)>>>(2'sd1)));

  assign y0 = ($unsigned((~|((&p9)?(b3):(3'sd3))))&((3'sd1)*((b0?b2:a0))));
  assign y1 = (|p9);
  assign y2 = ((a4?a3:a2)>>>(p0?a5:a2));
  assign y3 = (p9<p16);
  assign y4 = (((4'd4)-((p16<<<b0)!={b5})));
  assign y5 = {(5'd27),(-3'sd1)};
  assign y6 = {(({b4,b1,b0}===((a0|b0)|(a5+a1)))!==({(b4<b5),(a0>>>a4)}==={(b0<a5),(a4-b0)}))};
  assign y7 = (|(+(~&((+((p17&p17)<<((p6|p4))))))));
  assign y8 = (|(&({(({4{a3}}^(+b1))<<<((a1!=b4)+(p16<<a5)))}^{(({3{b2}}<<<(a2<<<b3))>=(-5'sd2))})));
  assign y9 = $signed(((((a3!==a4)>=(~p8))&&((a5-p11)||(a0-b0)))-$unsigned((!(((b2<=a5)&(p15^a0))-(!(-2'sd0)))))));
  assign y10 = ($unsigned({1{(p9==p13)}})||((a3===b5)+(b0==p13)));
  assign y11 = (((p3<a5)%p9)<((~((b0*b4)>>(5'd2 * b1)))>>((b4+b4)*(|p17))));
  assign y12 = {1{(-5'sd11)}};
  assign y13 = {1{((a1?a2:a0)?{2{a0}}:(p10^~b1))}};
  assign y14 = (b0?b2:b0);
  assign y15 = ((+(4'sd6))/b2);
  assign y16 = ({1{{p10,b5,p15}}}&({p1,p16,p16}==(-p17)));
  assign y17 = ((&{1{(~^(~^(!(!b4))))}})>{3{(p2?p5:p17)}});
endmodule
