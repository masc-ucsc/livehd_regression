module expression_00781(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(5'd1)}};
  localparam [4:0] p1 = {(-5'sd3),(3'd2),(-3'sd0)};
  localparam [5:0] p2 = ({((3'sd0)<<<(4'sd7)),((-5'sd12)<=(2'sd0))}<(4'd2 * ((2'd2)?(2'd2):(5'd2))));
  localparam signed [3:0] p3 = (((-4'sd0)>>((3'd6)<<(3'sd3)))^~((2'd0)<=(~|(-5'sd11))));
  localparam signed [4:0] p4 = (((-4'sd7)!=(3'sd0))^(!(-4'sd4)));
  localparam signed [5:0] p5 = {{(5'd13),(4'd6)}};
  localparam [3:0] p6 = {(4'd0),(-5'sd14)};
  localparam [4:0] p7 = ((((5'sd14)?(5'sd15):(-5'sd5))>>((3'sd3)==(2'd1)))<<(((2'sd0)/(3'd4))<<<((4'sd7)%(5'sd0))));
  localparam [5:0] p8 = {1{(4'sd1)}};
  localparam signed [3:0] p9 = (({2{(-2'sd1)}}|((-3'sd2)||(3'sd2)))!==(6'd2 * ((2'd1)?(3'd0):(5'd3))));
  localparam signed [4:0] p10 = {((4'd12)|(5'd8)),((-3'sd0)<=(3'd5)),(!(3'sd0))};
  localparam signed [5:0] p11 = (&((2'd1)===(-3'sd3)));
  localparam [3:0] p12 = ((3'sd3)!==(4'sd0));
  localparam [4:0] p13 = ({2{((-2'sd1)?(5'd18):(5'd3))}}?(!((4'sd5)?(5'sd1):(-5'sd14))):{2{((4'd12)&(3'd4))}});
  localparam [5:0] p14 = ({2{(5'd20)}}?((-4'sd7)?(5'sd5):(4'd12)):((5'd9)&(3'sd2)));
  localparam signed [3:0] p15 = {((3'd7)!==(3'd1)),((5'd9)<=(5'd11)),(6'd2 * (3'd5))};
  localparam signed [4:0] p16 = {1{{1{(~^{(^{((2'd2)<<<(-4'sd3))}),{1{(~&{(4'sd2)})}}})}}}};
  localparam signed [5:0] p17 = ((^(^(-4'sd3)))>(~&((-4'sd1)||(4'd9))));

  assign y0 = {(5'sd12)};
  assign y1 = (a3?p4:a0);
  assign y2 = (&(~&({(|a5),{a3,b4}}?(~&{a1,a2}):(~^{b4,b4}))));
  assign y3 = (2'd2);
  assign y4 = (~^((|$signed((&$signed((!p5)))))?((-(~(~^(p15?a5:p0))))):((~&b5)?$unsigned(p6):(p13?a3:a5))));
  assign y5 = ((^({{a2,a5,a3}}^~((-b3)===(~|a0))))<=(((b1==a3)&(a0+a0))||((a3&&a0)!==(4'd2 * b0))));
  assign y6 = (!(-((5'd12)?(3'sd3):(2'd1))));
  assign y7 = {(b4?b2:p1),(!b5),(a5?p1:a3)};
  assign y8 = (!((~&a3)?(|a5):{3{a5}}));
  assign y9 = {2{{(b0^a1),{{a2}},{p16,b4}}}};
  assign y10 = ((~($signed(((p8)?(p7?p2:b0):(p4<<<a1)))))+((3'sd2)?$signed((-2'sd1)):(-3'sd1)));
  assign y11 = (|(^(p9<<a0)));
  assign y12 = {(~|b1),{a5,p4,b0}};
  assign y13 = ((&(~&$unsigned((4'sd2)))));
  assign y14 = ((~^(~&(3'sd3)))?((~|a3)?(|p11):(3'sd0)):(4'sd4));
  assign y15 = (2'd0);
  assign y16 = ((b5?b3:b1)?({p4}<{b5,b3}):(a3?b0:p13));
  assign y17 = {(&p4),$unsigned(p3),(+b4)};
endmodule
