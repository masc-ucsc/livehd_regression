module expression_00786(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{((&(4'd2))>>((5'sd15)?(3'd0):(5'sd2)))}};
  localparam [4:0] p1 = (((&((4'sd3)&&(2'sd0)))>((-2'sd0)>>(5'd28)))<<<(((3'd1)>>>(3'd4))==((3'd6)^(2'sd0))));
  localparam [5:0] p2 = (({4{(3'sd2)}}!==((-2'sd0)<<(2'd0)))>=(~^(((4'd1)&&(-3'sd0))!=((5'sd11)>>>(-5'sd12)))));
  localparam signed [3:0] p3 = (|(((2'sd0)^(3'd3))<{(4'd0),(-3'sd2),(4'd11)}));
  localparam signed [4:0] p4 = ((|(2'd3))<<<(+(5'sd11)));
  localparam signed [5:0] p5 = (((((3'sd0)+(4'd1))||((3'sd1)^~(3'sd3)))>=(((4'sd7)==(4'sd1))^~((5'sd4)===(4'sd4))))^(((-4'sd2)|(3'd5))*((-4'sd1)+(4'sd5))));
  localparam [3:0] p6 = ((5'sd9)||(5'd28));
  localparam [4:0] p7 = ({(-(4'd0)),((2'sd1)<(-5'sd15)),((-3'sd0)>>>(4'd8))}|(~^{{(5'sd1),(5'd6)},{(2'd2),(5'd25),(-2'sd1)},((4'd11)<<(4'sd1))}));
  localparam [5:0] p8 = {1{(-2'sd0)}};
  localparam signed [3:0] p9 = (4'd15);
  localparam signed [4:0] p10 = (&((2'sd0)?(-5'sd2):(5'd15)));
  localparam signed [5:0] p11 = (-(6'd2 * (2'd3)));
  localparam [3:0] p12 = ((^(!((3'd1)?(5'd5):(-3'sd2))))?(~&((5'd12)<<(4'd8))):(~|(~|((5'd9)?(-5'sd14):(-3'sd2)))));
  localparam [4:0] p13 = ((-2'sd1)?(4'd0):(3'sd2));
  localparam [5:0] p14 = (4'd2 * ((5'd15)?(3'd7):(2'd0)));
  localparam signed [3:0] p15 = (-({1{(~{2{(-3'sd0)}})}}<<<(~&(~^((2'd3)!=(3'd3))))));
  localparam signed [4:0] p16 = {{1{((5'd9)^(5'd12))}},({3{(-4'sd0)}}+{(-2'sd0),(4'd13),(4'd4)}),{3{(-5'sd14)}}};
  localparam signed [5:0] p17 = (((-3'sd2)||((2'sd0)%(5'sd11)))>>(3'sd1));

  assign y0 = (|(~^(((~^a2)?(p17?p4:b1):(~^b2))?((b1||b1)?(~p4):(a5?a3:p5)):(~&(-(p12-a5))))));
  assign y1 = {(-(~p9)),(p12==a5)};
  assign y2 = (~(|((^(~|(&(a4*a4))))?$signed((a3?p5:a0)):(!(~&(b3^~a3))))));
  assign y3 = ((~&((((~|($signed((a5==b0))&(a2==b2))))>(((5'd2 * b0)|(a5-b4))&&{{(b2|a3)}})))));
  assign y4 = {(^({b3,a0,b3}?{b5,a0,b0}:{p1,a1,a4}))};
  assign y5 = (({a0,a0}==={a2,b4,a3})===({a3,a0}&(b4^~a5)));
  assign y6 = ((~^p3)<(p13-p1));
  assign y7 = (~&({(^(&(p12|p12)))}+((p10>>>p12)>(p3-p5))));
  assign y8 = {(b5?p5:b3),(p13||a1)};
  assign y9 = (+(~&(((&$unsigned($unsigned(p11)))<<<(~^(p14/p12)))|(!(&((5'd27)/p3))))));
  assign y10 = (a2?a4:a2);
  assign y11 = ((~&({b5,a1}?(a2!=a4):(p6?a0:a4)))<(((a2>>>a2))==(b2?b0:p11)));
  assign y12 = (|(5'sd8));
  assign y13 = ((5'd2 * $unsigned((~&a3)))^(+((^(a4>>b1))%b4)));
  assign y14 = (((&(^p0))*(^(b3^~p14))));
  assign y15 = {3{(&(3'd7))}};
  assign y16 = (2'sd1);
  assign y17 = (+{{({4{b1}}-(a2&p11)),({a2,b2}||(a4>=p8)),{2{(b0&p0)}}}});
endmodule
