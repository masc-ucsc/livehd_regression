module expression_00166(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+((3'sd3)?(-4'sd0):(3'd7)));
  localparam [4:0] p1 = ((~^(-4'sd4))>>>((5'd29)<=(4'sd6)));
  localparam [5:0] p2 = ((((2'sd0)!==(2'sd1))<{4{(3'd2)}})+({2{(4'd9)}}+((5'sd0)>=(-5'sd7))));
  localparam signed [3:0] p3 = (5'd26);
  localparam signed [4:0] p4 = ((-3'sd0)?(2'd3):(5'sd14));
  localparam signed [5:0] p5 = ((3'sd2)?(3'd5):(-4'sd0));
  localparam [3:0] p6 = ({4{(-3'sd1)}}|{4{(5'd20)}});
  localparam [4:0] p7 = (3'd2);
  localparam [5:0] p8 = {4{(5'sd3)}};
  localparam signed [3:0] p9 = (&(!((~((2'd1)<<(5'sd3)))?(|((4'd4)?(5'sd13):(4'd5))):((4'd15)?(-4'sd5):(4'd11)))));
  localparam signed [4:0] p10 = ((!(-5'sd3))<<(3'sd2));
  localparam signed [5:0] p11 = (~|(-2'sd1));
  localparam [3:0] p12 = {4{((2'sd0)^~(4'd7))}};
  localparam [4:0] p13 = ((+((-5'sd11)?(4'd11):(-4'sd3)))?(&(~(3'd7))):((5'd6)^~(4'd10)));
  localparam [5:0] p14 = {{(2'sd1),(2'd0)}};
  localparam signed [3:0] p15 = (-(-({3{(4'sd1)}}?{2{(5'd30)}}:{4{(2'sd1)}})));
  localparam signed [4:0] p16 = {(^(+(4'sd1)))};
  localparam signed [5:0] p17 = (&(-(~({(3'd4)}<<<((5'd0)<<<(4'd12))))));

  assign y0 = (p8&b0);
  assign y1 = (a0!==b4);
  assign y2 = (&(|((6'd2 * (p14>=a0))?(~(~|{a5,a3,b5})):(~^(b0?a4:b5)))));
  assign y3 = $signed((p9*p2));
  assign y4 = $unsigned((p11||a5));
  assign y5 = (!(-5'sd10));
  assign y6 = (|$unsigned((({4{a3}}?(+a2):(a3?p6:a4))&&(((~&b3)?(~a5):(+a1))))));
  assign y7 = (((|p8)==(~p15))<=((-3'sd2)<<<(-3'sd3)));
  assign y8 = ((&(^((!(p12%a3))>=((a5>p14)-(~p11)))))<<<((b0>b4)/b4));
  assign y9 = ((2'd0)<<(4'd2));
  assign y10 = ({4{a0}}<={3{{1{b4}}}});
  assign y11 = (((p16*a4)>>(a1^p2))|((p3*b0)>>>(~(a0+p6))));
  assign y12 = {(~^b4),(^b0),(&a3)};
  assign y13 = (3'sd0);
  assign y14 = ((3'd3)|{2{(4'd4)}});
  assign y15 = ({p5,p4,b1}?(b0?p13:p14):((a4===a4)+(a0||a4)));
  assign y16 = {{1{(a5!=p3)}}};
  assign y17 = ({2{p7}}>>(-4'sd7));
endmodule
