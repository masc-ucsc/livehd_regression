module expression_00137(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd0)?({(4'sd5),(5'd28),(5'd26)}>>>((-4'sd6)?(5'd26):(-3'sd3))):((5'd18)?(5'd6):(3'd5)));
  localparam [4:0] p1 = {({(-2'sd0)}-((4'd6)===(2'd3))),(((2'd1)>=(4'sd2))-{(3'd2)})};
  localparam [5:0] p2 = {(2'sd1),(-4'sd1),(3'd0)};
  localparam signed [3:0] p3 = (4'sd2);
  localparam signed [4:0] p4 = {1{(&(&{3{{2{(-3'sd2)}}}}))}};
  localparam signed [5:0] p5 = {4{(3'd6)}};
  localparam [3:0] p6 = (^((4'd12)?(-3'sd2):(!(-3'sd3))));
  localparam [4:0] p7 = (((5'd29)!=(5'd24))>=(!(2'd2)));
  localparam [5:0] p8 = ((-4'sd1)-(3'd0));
  localparam signed [3:0] p9 = ((-5'sd14)?(~^(4'sd7)):(!(2'sd0)));
  localparam signed [4:0] p10 = (-{{(~^{(3'd5),(2'sd1)}),((2'd0)&(-4'sd1))},((|((5'sd6)<(-3'sd0)))+{(2'd3),(3'd5),(4'sd6)})});
  localparam signed [5:0] p11 = {(3'd4),({(-5'sd8)}^~(5'sd5)),{{3{(2'sd0)}},{(-5'sd6)}}};
  localparam [3:0] p12 = {1{{{(4'd0),(-3'sd3),(5'd6)}}}};
  localparam [4:0] p13 = ((2'sd0)==(4'd2 * (4'd2)));
  localparam [5:0] p14 = ((~|(+(~^(-2'sd1))))?(&(-((3'd1)<=(3'sd0)))):((&(5'sd15))<(~(5'd5))));
  localparam signed [3:0] p15 = ((~{(&{(4'sd7),(2'sd0),(4'd0)})})!==(|((+(4'sd6))>>{(4'd1),(2'sd0),(4'd4)})));
  localparam signed [4:0] p16 = (~|(5'sd1));
  localparam signed [5:0] p17 = ((&(~|{2{(|{1{(3'd1)}})}}))<<(|{2{((5'd20)^(4'd10))}}));

  assign y0 = (~|(-2'sd0));
  assign y1 = {3{{(b2^b5)}}};
  assign y2 = (4'd2 * (b1^~b2));
  assign y3 = (($signed($unsigned((a0|a4)))!={(a1<a5),{b0,a4}}));
  assign y4 = {(-{4{p2}}),(!(&(-p8)))};
  assign y5 = (p9>p1);
  assign y6 = ($signed(((|(a4<a0))/a5))+$unsigned((+(-$unsigned((~((+p9))))))));
  assign y7 = (~|(^{2{{2{{3{b4}}}}}}));
  assign y8 = {$unsigned((-{b4,a0,a1})),{(a0>>b2)}};
  assign y9 = (((&(a1<=b3))<<<(b2!==b5))>=(~&{2{{4{a2}}}}));
  assign y10 = ((-5'sd6)?(3'sd0):(b4>a4));
  assign y11 = {2{((a5?p13:p5)?{3{p8}}:(p3+a1))}};
  assign y12 = ((a3||a3)+(b5>>b5));
  assign y13 = (2'd1);
  assign y14 = ((~^(3'd2))>>(((-5'sd0)>>>(+b4))>>>((2'd2)!==(4'd8))));
  assign y15 = (((a0!==b5)%p12)?(-((p7<=p15)^(p15/p2))):((p11/p13)%p7));
  assign y16 = {(((+a5)>{b2,b1,b4})>>((~|b3)<<<(^b2))),(((a2<<b3)<={3{b2}})|({a1,b4}-{3{b4}}))};
  assign y17 = ({4{$signed($unsigned({a4}))}});
endmodule
