module expression_00353(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-5'sd9);
  localparam [4:0] p1 = ((2'd0)==(2'sd0));
  localparam [5:0] p2 = ((3'd6)<=(4'd8));
  localparam signed [3:0] p3 = ((4'd6)!=(4'd6));
  localparam signed [4:0] p4 = {3{((5'd9)?(4'd5):(5'd17))}};
  localparam signed [5:0] p5 = ((~|(3'd5))+((-5'sd12)==(3'd0)));
  localparam [3:0] p6 = (((5'd20)>>(3'd1))>=(3'sd0));
  localparam [4:0] p7 = (((6'd2 * (4'd14))>>>(+(5'd22)))===(5'd2 * ((3'd6)&(5'd28))));
  localparam [5:0] p8 = ((6'd2 * (4'd12))==((2'sd0)<(5'sd6)));
  localparam signed [3:0] p9 = {(2'd3),(4'd12)};
  localparam signed [4:0] p10 = (2'd3);
  localparam signed [5:0] p11 = (+(2'd3));
  localparam [3:0] p12 = (+({(^(~|(+(-3'sd1))))}==(|{(5'd31),(-2'sd0),(5'd2)})));
  localparam [4:0] p13 = (~&(!(|(~(~|(+(5'sd8)))))));
  localparam [5:0] p14 = ((5'd8)==(5'sd9));
  localparam signed [3:0] p15 = {{{(-4'sd1)},{(3'd4),(-3'sd0),(3'sd3)}}};
  localparam signed [4:0] p16 = (((-5'sd6)?(4'sd6):(2'sd0))?{2{(-5'sd9)}}:{2{(5'd17)}});
  localparam signed [5:0] p17 = {1{{1{(-(2'd2))}}}};

  assign y0 = (~({4{(-4'sd1)}}||(5'd2)));
  assign y1 = {{(2'd2)},($signed(a0)-(4'sd7)),((p11!=p2)!=(p2|a0))};
  assign y2 = (a1?p2:b3);
  assign y3 = (((b0)%p14)?((b3-b5)):(~^(b2<<<b0)));
  assign y4 = (p4&a3);
  assign y5 = ({(!(p7==p10)),{p1,p9},(p6<p1)}<<<{(-((p12?p3:p8))),$unsigned((p13!=p1))});
  assign y6 = (^({{3{p11}},(p8||p8)}?(&(!(-(!p5)))):{{2{p17}},(!p17),(p17>=p16)}));
  assign y7 = {4{(b2!=a4)}};
  assign y8 = (~^({3{(~&a1)}}?{2{(^(~^p3))}}:(-2'sd1)));
  assign y9 = (((4'sd3)?(p0*p3):(p7?p7:a3))?(2'd0):((b5?p6:p13)?(-3'sd2):(b3?b4:a2)));
  assign y10 = ({b4,b0,a1}==={4{b2}});
  assign y11 = (~^(^(3'd6)));
  assign y12 = ((~|(-2'sd1))^(~|(-3'sd3)));
  assign y13 = $unsigned((3'sd1));
  assign y14 = {1{{2{(5'sd4)}}}};
  assign y15 = ({3{p13}}?{4{p2}}:$signed(a1));
  assign y16 = (p5);
  assign y17 = {2{{3{$unsigned({3{a1}})}}}};
endmodule
