module expression_00335(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd5)+(2'sd1));
  localparam [4:0] p1 = (((2'd0)<<<(2'd3))===((5'd19)<<<(5'd20)));
  localparam [5:0] p2 = (-{4{(|{1{(-2'sd0)}})}});
  localparam signed [3:0] p3 = (2'd1);
  localparam signed [4:0] p4 = {2{(((4'd5)|(4'd7))?((4'sd2)>>(3'sd2)):{4{(-3'sd0)}})}};
  localparam signed [5:0] p5 = ((3'sd3)&&(((2'd1)<<(5'd15))==={2{(2'd2)}}));
  localparam [3:0] p6 = (((&((2'd0)-(4'd0)))+(~(~(5'd1))))&&((^(-2'sd1))?{3{(-5'sd1)}}:(~(2'd0))));
  localparam [4:0] p7 = (^(2'd0));
  localparam [5:0] p8 = (~^(^(|(~(~((4'd3)|(-3'sd2)))))));
  localparam signed [3:0] p9 = {{((-3'sd2)!=(5'd7)),((4'd5)?(4'd7):(5'd5)),((5'd5)?(3'd7):(5'sd12))}};
  localparam signed [4:0] p10 = (~^(&(!(4'sd1))));
  localparam signed [5:0] p11 = ((5'sd8)===(3'd1));
  localparam [3:0] p12 = {((2'd2)+(5'd24)),((4'd3)<=(3'sd0)),((5'd25)^(5'd6))};
  localparam [4:0] p13 = {{(&(2'd3)),((4'sd6)<=(2'd3))},(~|(~&{(-5'sd10),(5'd13),(2'd3)})),((~(3'sd0))!==(~|(5'd1)))};
  localparam [5:0] p14 = (3'sd2);
  localparam signed [3:0] p15 = ((4'sd3)===(5'sd4));
  localparam signed [4:0] p16 = {3{(((-5'sd5)>>>(5'd3))<<((2'd1)||(2'sd1)))}};
  localparam signed [5:0] p17 = ({3{(-2'sd0)}}+{2{(-4'sd3)}});

  assign y0 = {1{(~&(&p10))}};
  assign y1 = (b4<<b5);
  assign y2 = {1{{2{((a1>>a4)^{a5,a5,b3})}}}};
  assign y3 = ((~|(|(~(&(3'd1)))))<(2'sd0));
  assign y4 = {1{(({1{b0}}==(b4<<b4))?((b4===a3)+{a3}):({a3}>>(b1?b4:a0)))}};
  assign y5 = ({$signed(p2),(a3!==b3)}?((p7==p11)<<(p10?p2:p13)):(p10?p3:p1));
  assign y6 = ($unsigned({4{$signed(a4)}})-(({4{p2}}=={4{a3}})!=({4{a5}}>=(~^b5))));
  assign y7 = (~|(-(p11?p1:p0)));
  assign y8 = {{2{{4{p15}}}},{4{{a5,a5}}}};
  assign y9 = (((a4>>a0)&&(p4!=p6))|((b1|a2)%a4));
  assign y10 = ((((4'd2 * a0)&&(a4&&a4))>((b5===b0)!==(a3|a3)))!==(((a2||b0)&&(b5+b1))<<((a5<<b1)|(b3&&b5))));
  assign y11 = {(&(p10?p1:p1)),({p4,p0}?(-p9):(p2?p4:p12))};
  assign y12 = (!{((p15>p5)+(p4||b4)),{(p3>>>p7)},$signed({p4,p1,p10})});
  assign y13 = (((p3)?(!p7):(b0?b5:p0))?((-((2'd2)-$signed(a0)))):((-5'sd5)?(&a5):(2'd1)));
  assign y14 = {4{(2'd2)}};
  assign y15 = (+(&b3));
  assign y16 = (~|(((2'd2)?(~&b5):(3'd5))-((b0?a4:b3)?(a3?a4:b2):(a0+b0))));
  assign y17 = {2{{{a5,p10},$unsigned(a2)}}};
endmodule
