module expression_00647(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|((!(|{(~^(-(-3'sd0)))}))&&(~&((|(4'd15))-(~&(4'd3))))));
  localparam [4:0] p1 = {(-5'sd2),(-2'sd1),(-5'sd6)};
  localparam [5:0] p2 = ((~(~|(((2'd3)!=(-4'sd2))+(~^{1{(-4'sd6)}}))))|(((~&(2'sd0))<={1{(5'd9)}})===(!{4{(2'd3)}})));
  localparam signed [3:0] p3 = ((&((-2'sd0)?(-4'sd0):(-5'sd9)))===({2{(-5'sd9)}}?{4{(4'd15)}}:(~^(-4'sd2))));
  localparam signed [4:0] p4 = (-5'sd8);
  localparam signed [5:0] p5 = (~|((((-3'sd0)>>(2'sd1))<<<{(-5'sd4),(4'sd6),(5'd21)})<=(((2'sd1)?(2'd0):(-3'sd1))||((3'sd2)?(-2'sd0):(2'd0)))));
  localparam [3:0] p6 = {1{(4'd2 * {(3'd2),(2'd0)})}};
  localparam [4:0] p7 = {3{(3'd6)}};
  localparam [5:0] p8 = (((-2'sd0)<=(5'd1))/(5'd17));
  localparam signed [3:0] p9 = ((4'd1)?{(5'd5),(5'sd11),(3'd4)}:{{(5'sd11),(4'd15),(3'sd0)}});
  localparam signed [4:0] p10 = ((4'd6)>>>((|(-4'sd1))==((3'd2)-(2'd0))));
  localparam signed [5:0] p11 = {(3'd7),(2'd1)};
  localparam [3:0] p12 = (((3'sd1)?(3'sd0):(-2'sd0))?((4'sd0)?(-4'sd7):(3'sd0)):((3'd4)?(2'sd1):(-5'sd1)));
  localparam [4:0] p13 = (-5'sd6);
  localparam [5:0] p14 = (~&((~|((5'd24)%(3'd4)))^((&(-2'sd0))+(~&(3'd5)))));
  localparam signed [3:0] p15 = {{(2'sd1),(3'd2),(4'sd4)},{(3'sd2),(4'sd2),(-2'sd0)}};
  localparam signed [4:0] p16 = (2'd1);
  localparam signed [5:0] p17 = (((~^((2'd1)?(4'sd3):(-5'sd2)))*(&(3'sd0)))!==(((4'd5)<=(5'd8))<(3'd0)));

  assign y0 = {3{{3{{4{p6}}}}}};
  assign y1 = ((-4'sd1)||(3'sd2));
  assign y2 = (5'sd4);
  assign y3 = (((b3||p10)&{p13,a4})>>>(((a0&p14))<={p16,a1,b4}));
  assign y4 = (^(((b1?p3:p2)?(4'd13):(b0?p0:p1))&(3'd1)));
  assign y5 = ((p4?p8:p3)?(p17>b2):(b0|a5));
  assign y6 = (((5'd2 * (a1>>a0))>(~^{(b2>>>a4),(&b2),$signed(a3)})));
  assign y7 = ((((p3>=b5)-(b5^~a1))!=((p14>=a3)/p15))+(((b0!=p5)%b2)&&((b4&b5)>=(p16<<<a1))));
  assign y8 = (4'd14);
  assign y9 = {3{(&({3{p5}}+{1{{p9,p13,p17}}}))}};
  assign y10 = (+(^(~&(&(3'd4)))));
  assign y11 = (({b0,b1}?(6'd2 * a2):(-a5))-((p5?p9:b0)-(p12^b3)));
  assign y12 = ({1{{(a3===a0),(a2||a1)}}}-(-{(a3?a1:a3)}));
  assign y13 = ((~&((b5?b5:b2)===(&(a1+b0))))?(~{(~((b3?b5:a5)^{a0}))}):((a5?b2:b1)<={a4,b4,a0}));
  assign y14 = (5'd22);
  assign y15 = {1{(~((p0>=p8)<<(~&(a3===b0))))}};
  assign y16 = (3'd7);
  assign y17 = ($signed({(-$signed($signed(a1)))})?($unsigned((~|(b1?a4:a1)))):$unsigned({{b0,b3},(b2)}));
endmodule
