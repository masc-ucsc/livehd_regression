module expression_00350(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd5);
  localparam [4:0] p1 = (5'sd6);
  localparam [5:0] p2 = (~&((((5'sd1)-(5'd13))?{1{(-5'sd1)}}:{1{(5'd22)}})?(3'sd1):({4{(4'd10)}}?{3{(4'sd3)}}:{1{(3'sd3)}})));
  localparam signed [3:0] p3 = (5'd25);
  localparam signed [4:0] p4 = (|(~^(~(~(5'd29)))));
  localparam signed [5:0] p5 = ((5'd18)?(2'sd1):(-5'sd12));
  localparam [3:0] p6 = {{{(-2'sd0),(4'd15)}},{2{(4'sd5)}}};
  localparam [4:0] p7 = (~&(+(~(+(~|((-{(-5'sd8)})!=((-3'sd0)===(5'd8))))))));
  localparam [5:0] p8 = (&((-(-2'sd0))?(^(4'd9)):(2'sd0)));
  localparam signed [3:0] p9 = (+{1{(4'd3)}});
  localparam signed [4:0] p10 = {(5'sd2)};
  localparam signed [5:0] p11 = (~(2'd0));
  localparam [3:0] p12 = ((4'sd0)?(4'sd0):(-3'sd3));
  localparam [4:0] p13 = ((4'd4)<={((4'd4)|(-3'sd3)),(-(-5'sd10))});
  localparam [5:0] p14 = ((-(~&(-3'sd0)))?((-5'sd0)?(2'sd0):(5'd1)):((2'd3)?(3'sd0):(3'sd1)));
  localparam signed [3:0] p15 = (^({1{((~&(2'd3))<{1{(2'sd1)}})}}<=((&((4'd12)>=(2'sd0)))-{3{(4'sd0)}})));
  localparam signed [4:0] p16 = (((~|(5'd30))<<<(~(-3'sd1)))<<<((|(3'sd2))<((-4'sd5)==(5'd17))));
  localparam signed [5:0] p17 = (({4{(-4'sd5)}}<{4{(4'd9)}})<<<{2{{3{(2'd1)}}}});

  assign y0 = ((~^{{4{p14}}})^({1{{b0}}}|(+{p5,p9,p13})));
  assign y1 = ((b1==a3)|(p14?b1:b2));
  assign y2 = (3'd1);
  assign y3 = $unsigned({{(p10-p17),(p1^~p13)},{{p14,p5},(~p13),{p10,p13}},{(-(p2)),(p13?p15:p7)}});
  assign y4 = (($signed((a5&b4))));
  assign y5 = (4'd14);
  assign y6 = ((5'd18)>=(((p10*p9)-(b4?b4:b4))&((p13?a5:p1)<<<(p6-b5))));
  assign y7 = {b2,a1};
  assign y8 = ((5'd24)<=(p6?p5:p15));
  assign y9 = ((p8&&p9)<={p16,p15});
  assign y10 = (-(+(((~|p0)<<<(!a2))?(~(p7<=a0)):(~(p16?p3:p10)))));
  assign y11 = ((5'd2 * {b0,p2})!=({{p5,b1}}>>$unsigned((~^(p17^a3)))));
  assign y12 = {p3,p2};
  assign y13 = (2'd2);
  assign y14 = {3{(-2'sd0)}};
  assign y15 = (&{2{a1}});
  assign y16 = ((^$unsigned($signed((p7))))<<<(+(p16?b3:a1)));
  assign y17 = $signed({{$signed(p15),{3{p8}}}});
endmodule
