module expression_00816(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-4'sd2)?(-2'sd0):(3'd6))?(5'd27):(3'd6))<<((5'd5)===((5'd24)^~(-2'sd1))));
  localparam [4:0] p1 = (^(4'd11));
  localparam [5:0] p2 = (2'sd0);
  localparam signed [3:0] p3 = {(|((3'd0)&(-3'sd3))),(((5'd8)^~(5'd16))>=((3'sd1)>>(-3'sd1))),(+{(4'd0),(-4'sd6),(-5'sd12)})};
  localparam signed [4:0] p4 = ({4{((3'sd1)?(2'd2):(5'sd3))}}<<<(((5'd4)>(2'd0))?((-4'sd5)?(3'd4):(2'sd0)):((-2'sd1)?(-3'sd1):(3'd7))));
  localparam signed [5:0] p5 = (({(-4'sd3),(4'd14)}<(&((4'd2)>>>(3'd0))))==({((-2'sd0)||(3'd7))}+(4'd4)));
  localparam [3:0] p6 = (^(-3'sd0));
  localparam [4:0] p7 = ({(+{(4'sd3),(-3'sd1)})}>>{4{(-2'sd1)}});
  localparam [5:0] p8 = (!(5'sd10));
  localparam signed [3:0] p9 = ({3{(5'd15)}}?((-3'sd0)|(3'sd2)):((2'sd1)<<(-4'sd2)));
  localparam signed [4:0] p10 = ((~((-4'sd6)?(2'd1):(4'sd2)))?((2'd0)?((-3'sd0)?(5'd22):(-5'sd0)):(~(3'd5))):((~^(-5'sd1))!=((-5'sd7)==(2'sd0))));
  localparam signed [5:0] p11 = ((2'd2)?(2'd1):(3'd2));
  localparam [3:0] p12 = (3'sd3);
  localparam [4:0] p13 = (((4'sd7)^(-2'sd1))>(4'd2 * (3'd1)));
  localparam [5:0] p14 = (&(((+((3'sd1)!=(-2'sd0)))^((-4'sd7)>>(5'd19)))===((-((4'd13)!=(2'd1)))&&(~^((5'sd11)*(-2'sd0))))));
  localparam signed [3:0] p15 = ({(2'd2),(-4'sd3),(-4'sd3)}!={((5'd2)|(-2'sd1))});
  localparam signed [4:0] p16 = (~^({(-(-4'sd3)),((3'd1)?(-2'sd0):(3'd2))}?((^(4'sd7))?((-4'sd7)?(2'd2):(5'd0)):{(-2'sd0),(2'sd0)}):(-(~|{(5'sd0),(2'd0)}))));
  localparam signed [5:0] p17 = {1{(-{2{(~(-(3'sd2)))}})}};

  assign y0 = ((4'd2 * {3{b1}})>>(2'sd0));
  assign y1 = ($signed((4'd2 * b2))*(!(-a4)));
  assign y2 = ({b3,b5,a1}==={4{a4}});
  assign y3 = (~|(~&(~|({1{{1{((a5<<<p13)^{4{p5}})}}}}!=(|(~|((|(b1&&a0))<<<(~|(p12>>p14)))))))));
  assign y4 = (|{p17,b0,p2});
  assign y5 = ((~&{2{(~&p14)}})-({1{p11}}&(p4^~p3)));
  assign y6 = (((b0-p5)<<(~|a4))>=((p9^b3)-(a1<=a1)));
  assign y7 = (4'd12);
  assign y8 = ((p17&&p10)?(a5===b3):(b5?p1:b2));
  assign y9 = {{(5'd31),((p8||p2)>(-4'sd3))},(-4'sd0)};
  assign y10 = {({2{b4}}<={1{p17}}),{4{p0}}};
  assign y11 = $signed(($signed($unsigned((~&((p11?b4:p10)?(~(b0?b5:p8)):((b0<p10)-(p3?a3:a2))))))));
  assign y12 = {1{(($signed({p13,p1}))==((2'd0)>>{p0}))}};
  assign y13 = $unsigned(((p1?p0:p5)?((&(p2?p11:p7))):(p10?p5:p1)));
  assign y14 = (|(-2'sd1));
  assign y15 = (p3?a5:p15);
  assign y16 = {4{p1}};
  assign y17 = {2{(^{b2,p13,b2})}};
endmodule
