module expression_00242(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((5'sd1)<<<(5'd19))|((-5'sd10)<=(-5'sd15)))-({(2'd1),(4'd5)}!={(4'd12)}));
  localparam [4:0] p1 = (~|((4'd4)>={4{(-4'sd2)}}));
  localparam [5:0] p2 = (-((|(5'd20))>=(-2'sd1)));
  localparam signed [3:0] p3 = (!((5'd23)?(-3'sd2):(-3'sd3)));
  localparam signed [4:0] p4 = (~&{(5'd2 * ((4'd11)?(4'd5):(2'd0)))});
  localparam signed [5:0] p5 = (3'sd0);
  localparam [3:0] p6 = (5'd2 * (5'd10));
  localparam [4:0] p7 = (+(-3'sd1));
  localparam [5:0] p8 = (6'd2 * ((2'd3)>>>(3'd2)));
  localparam signed [3:0] p9 = (|((+(&(~&(^((-2'sd0)||(3'd2))))))>>>({2{(2'd1)}}^((5'd4)^~(-5'sd9)))));
  localparam signed [4:0] p10 = (4'd5);
  localparam signed [5:0] p11 = (-(5'd24));
  localparam [3:0] p12 = (4'sd3);
  localparam [4:0] p13 = (3'd2);
  localparam [5:0] p14 = ((&(~(((2'd1)===(-2'sd0))?(~^(-3'sd2)):(~&(4'd10)))))^~(^(((5'sd0)>=(4'sd1))&(-(~^(3'sd0))))));
  localparam signed [3:0] p15 = {3{(+{2{{1{(3'd5)}}}})}};
  localparam signed [4:0] p16 = (((3'd3)>(3'd6))===(+((5'd16)<(5'sd6))));
  localparam signed [5:0] p17 = ((4'd9)?(5'sd6):(2'd0));

  assign y0 = (+((-2'sd0)?(5'sd1):(p11?p11:p13)));
  assign y1 = ($unsigned((+(b0==p5)))^$unsigned((p15-p4)));
  assign y2 = (2'sd1);
  assign y3 = (~^(~|(!((~^(($unsigned($unsigned(b1))>>$unsigned($signed(b4)))!==(((a5===a3))==$signed((a2|a3)))))))));
  assign y4 = ((b0?a3:a4)>=({b1,b5}<(2'd1)));
  assign y5 = (&(^{(!(-4'sd2))}));
  assign y6 = (((p13==p12)&&(a0<<p9))>((p13^b4)^(p3<<<p14)));
  assign y7 = {1{(((6'd2 * a0)==(-b5))!==(-2'sd1))}};
  assign y8 = (~&((|({b4,b5,b0}&(5'sd3)))+(4'd15)));
  assign y9 = ((a5+a4)&(b3<b2));
  assign y10 = (b1/b3);
  assign y11 = (a0?b4:b2);
  assign y12 = ({{3{{1{p9}}}},((a2)^~(p10))}&{1{(~{1{{4{{p7,a0}}}}})}});
  assign y13 = {b3,p17};
  assign y14 = (~^((!{a4,a2,p12})^({2{p4}}>>>{4{p5}})));
  assign y15 = (|(({a4,p10,p12}|((b2!==a1)!=(b5!==a4)))<={{(^b4),(p16<<p0)},$signed({p14,p9})}));
  assign y16 = (((b5>a5)<<<{4{a3}})!==$unsigned((b1<=b5)));
  assign y17 = (((b3!==a0)+(a4>p1))>>((a2>>p7)>(~a3)));
endmodule
