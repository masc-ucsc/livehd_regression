module expression_00429(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~(+{2{(-3'sd0)}}))-((5'sd15)?(5'd10):(2'sd0)));
  localparam [4:0] p1 = {4{(~^(|(-4'sd1)))}};
  localparam [5:0] p2 = ((4'd2)>>((&(5'sd14))-((-3'sd1)-(-3'sd0))));
  localparam signed [3:0] p3 = (({4{(5'sd11)}}|((3'd7)<=(3'd6)))>>>(((5'sd5)?(5'sd11):(5'd8))<(5'sd2)));
  localparam signed [4:0] p4 = (~(({2{(5'd23)}}^{2{(2'd3)}})?{2{{3{(-4'sd2)}}}}:(|(&((2'd0)<=(3'sd2))))));
  localparam signed [5:0] p5 = {4{{4{(5'd26)}}}};
  localparam [3:0] p6 = ((~|{2{(-5'sd9)}})=={(3'd3),(5'd7),(5'd14)});
  localparam [4:0] p7 = (&(&(~&(-(+(-(+(+(3'sd3)))))))));
  localparam [5:0] p8 = (~|(~^(6'd2 * ((4'd5)<=(3'd3)))));
  localparam signed [3:0] p9 = ((3'd5)<<(3'd7));
  localparam signed [4:0] p10 = {4{(3'd5)}};
  localparam signed [5:0] p11 = (4'sd2);
  localparam [3:0] p12 = (~(((!(5'd17))==(+(-5'sd8)))!==(+((-2'sd0)!==(5'd14)))));
  localparam [4:0] p13 = ({2{(2'd1)}}>((3'sd1)?(4'sd4):(3'd0)));
  localparam [5:0] p14 = ((5'sd8)?{2{{(4'd0),(5'd25),(2'd3)}}}:{((-2'sd1)?(2'sd0):(-5'sd5))});
  localparam signed [3:0] p15 = {{(((3'sd2)&&(4'sd5))?{(-2'sd0),(3'sd2)}:(~^(4'd10))),((5'd2 * (3'd1))?{(-4'sd6)}:((3'd0)+(5'd11))),(((-2'sd0)>>(3'd3))=={(2'd0),(4'd2)})}};
  localparam signed [4:0] p16 = {(&(2'sd0)),((2'd0)||(5'd1)),(5'sd13)};
  localparam signed [5:0] p17 = ({(4'd11),(5'd1),(3'sd2)}<((3'sd0)>>(3'd1)));

  assign y0 = (4'd9);
  assign y1 = ({(+a2),{1{a3}},(|p1)}?((b2>p3)&{p12,a5}):((a5^p14)!=(|{p5,b2})));
  assign y2 = (&(5'd16));
  assign y3 = ({{(-{(!(&a3))}),(-(~^(~|(|p13)))),{(^$signed({p2,a5}))}}});
  assign y4 = ((2'd1)!==(+a1));
  assign y5 = ((b5?a4:a1)?((2'sd0)>>(4'sd1)):((2'sd0)|(3'sd2)));
  assign y6 = (-(|(+(2'd1))));
  assign y7 = {1{{1{(4'd5)}}}};
  assign y8 = ({a4,b3}<$unsigned(a0));
  assign y9 = ((-(~|(~&((~|$unsigned((b3)))!==((b5||b3)>={4{a4}}))))));
  assign y10 = ((((^b0)||(a1<b1))<(-2'sd1))!=(-(((5'd4)|(a4^~a0))===(3'd2))));
  assign y11 = {{a2,b2,b5},{2{a3}},(3'd6)};
  assign y12 = {1{$unsigned({4{(3'sd3)}})}};
  assign y13 = (+(5'd2 * (b2-p8)));
  assign y14 = (p12?a4:a3);
  assign y15 = ($signed((p13)));
  assign y16 = $signed({4{($signed(b3)?(b2>>>a4):{4{b3}})}});
  assign y17 = (2'sd0);
endmodule
