module expression_00256(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^((4'd9)+(4'sd5)))<<<(((4'd15)===(3'sd3))&&(5'd7)));
  localparam [4:0] p1 = (((3'd6)?(5'd10):(4'd9))<((5'd11)?(4'd9):(-5'sd7)));
  localparam [5:0] p2 = {(5'sd9)};
  localparam signed [3:0] p3 = (((-5'sd9)<<<(5'd6))?((4'd14)-(2'd2)):{(5'd2),(3'sd1)});
  localparam signed [4:0] p4 = (5'sd7);
  localparam signed [5:0] p5 = {{2{{2{{2{(4'd3)}}}}}}};
  localparam [3:0] p6 = {((&{(3'd2),(3'd1),(5'sd7)})^~{{(-4'sd3),(4'sd1)}}),(|(^{(+((5'd21)>=(-5'sd8)))}))};
  localparam [4:0] p7 = (({4{(2'sd0)}}>=(!(3'sd1)))+(|((5'd5)>=(-3'sd2))));
  localparam [5:0] p8 = (-2'sd1);
  localparam signed [3:0] p9 = (-4'sd5);
  localparam signed [4:0] p10 = (~^(2'd2));
  localparam signed [5:0] p11 = (-3'sd2);
  localparam [3:0] p12 = (((3'd2)^(-2'sd0))%(5'd2));
  localparam [4:0] p13 = (((2'sd1)-(-3'sd1))<<<((5'sd14)?(4'd6):(5'd18)));
  localparam [5:0] p14 = (-5'sd4);
  localparam signed [3:0] p15 = (({(5'sd4)}|((3'sd2)==(4'sd5)))<(((3'sd2)+(-2'sd0))<{(5'd29),(3'd7)}));
  localparam signed [4:0] p16 = {(3'sd3)};
  localparam signed [5:0] p17 = (~&{(-5'sd8),(2'd2)});

  assign y0 = (|(-(~&a4)));
  assign y1 = ((p17&&b1)?(p2^p15):(b4===b5));
  assign y2 = ($unsigned((6'd2 * p14))>(-(a3===a2)));
  assign y3 = ({((b0|a4)<(b3!==a0)),(p2?a2:b3)}==((a3!==a0)?(a4===a0):{(b3-a5)}));
  assign y4 = $signed({4{$signed(b5)}});
  assign y5 = ((5'sd2)>{p15,b1,p3});
  assign y6 = ($signed(($unsigned(((b4?a4:b5)?$unsigned(p12):(p3?p16:b1)))?((a4?a1:b5)?(b4?p3:p15):(p11?a3:a3)):((p1?p10:p7)?$unsigned(p11):(p10?a0:b0)))));
  assign y7 = ({1{a2}}^~{2{p11}});
  assign y8 = {3{{3{(p17?a0:p0)}}}};
  assign y9 = (-4'sd0);
  assign y10 = (~^{4{(p9?b4:p6)}});
  assign y11 = ((-3'sd3)?((b2?b2:a2)<<(|p8)):(-((~^p2)<<(-3'sd2))));
  assign y12 = (b3<b3);
  assign y13 = {2{{1{(+(p12>>p3))}}}};
  assign y14 = ((5'd2 * p0)<<$signed($unsigned(b1)));
  assign y15 = (3'd4);
  assign y16 = $signed((^(-4'sd7)));
  assign y17 = (!(4'sd0));
endmodule
