module expression_00223(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((^(4'sd2))?{{(2'sd1),(2'd0),(4'sd2)}}:(2'sd1))=={((~^(-2'sd0))<<<((3'sd2)?(4'sd0):(-4'sd0))),{((5'd22)==(4'd2))}});
  localparam [4:0] p1 = {3{(&(|(+{2{(4'd10)}})))}};
  localparam [5:0] p2 = {({(4'sd4)}^~((4'd15)^~(4'd3))),(|((2'd2)!==(5'd25)))};
  localparam signed [3:0] p3 = {2{{{3{(2'd2)}},{3{(4'd2)}},{(-2'sd0),(4'sd1),(2'd2)}}}};
  localparam signed [4:0] p4 = (~^(((4'd6)^(4'sd2))||((4'sd0)>=(-4'sd6))));
  localparam signed [5:0] p5 = {(5'd16)};
  localparam [3:0] p6 = {(~|(-{((-(3'sd3))^~(&(2'sd1))),(|(~{(-3'sd0)})),((~|(2'd3))<((4'd7)<=(5'sd2)))}))};
  localparam [4:0] p7 = (4'sd4);
  localparam [5:0] p8 = (~^(^(-5'sd13)));
  localparam signed [3:0] p9 = (!(~|((3'd7)?(4'd4):(2'sd1))));
  localparam signed [4:0] p10 = (5'sd10);
  localparam signed [5:0] p11 = (6'd2 * (5'd2));
  localparam [3:0] p12 = {{4{{((3'sd3)?(-2'sd1):(3'd0)),((5'd1)>(-5'sd0))}}}};
  localparam [4:0] p13 = (((5'd13)!=={(4'sd4),(-5'sd13),(5'd16)})>=((2'sd0)-{(3'd0),(-3'sd1),(4'sd4)}));
  localparam [5:0] p14 = (!({((-4'sd6)<<<(5'd27)),(&(-2'sd1)),(!(4'd10))}^({(3'd7),(-5'sd8)}^{1{((-5'sd12)<<<(3'd4))}})));
  localparam signed [3:0] p15 = {(+((3'd4)<(2'sd1)))};
  localparam signed [4:0] p16 = {(({(3'd4)}==(~|(-4'sd6)))===(((-2'sd0)|(3'sd2))^{(-5'sd1),(2'sd0)}))};
  localparam signed [5:0] p17 = ((~&(((-5'sd5)==(5'd13))!=={(4'd2),(2'd2)}))|(4'sd0));

  assign y0 = (|({1{((|((a3?a5:a4)?(b5<<a3):(b1<a3)))^(~^{4{(b2>>>b1)}}))}}));
  assign y1 = {((^$signed((+(-$signed($signed(((-$unsigned((~^(^(+$unsigned((~^(!p15))))))))))))))))};
  assign y2 = (!(~|((~^($unsigned(p5)?{2{p3}}:(!p16)))?$signed(($signed(p7)?(p14):(b3===a0))):((~|(p10?p9:p2))!=(p10?p11:p4)))));
  assign y3 = (!(((a5===b2)||$unsigned(p2))^{4{p9}}));
  assign y4 = {b5};
  assign y5 = {{(~&((~^p13)^~{p15,p12}))}};
  assign y6 = ((2'd2)||{4{(5'd10)}});
  assign y7 = {2{{{3{(b3==p15)}},(~({b5,b5,b1}==(p10-p11)))}}};
  assign y8 = ((b0?b2:b3)?(a2?b3:a1):(b3?a2:b5));
  assign y9 = ((p16^~a4)<(p9^~b3));
  assign y10 = {3{{2{b5}}}};
  assign y11 = (3'd4);
  assign y12 = ((-5'sd0)?{3{b5}}:(a3?b2:p3));
  assign y13 = {($signed((b5>>>a0))?(b2>>>b1):(b5<b0))};
  assign y14 = (2'd0);
  assign y15 = $unsigned(p13);
  assign y16 = {((p16^~b3)+$signed((p8+p5))),(4'd5),{(!{{p15,p11,p16}})}};
  assign y17 = (^(!(!(~(~(&(+(^(|(!p14))))))))));
endmodule
