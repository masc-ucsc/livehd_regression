module expression_00827(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'd7)-(-2'sd1))==((2'd2)|(3'sd3)));
  localparam [4:0] p1 = (((5'd2)!==(2'd0))*((5'd4)?(5'sd14):(5'd20)));
  localparam [5:0] p2 = (~&((~&(~{4{(5'd0)}}))|(|((4'sd1)&&(~((3'd1)?(4'd7):(-3'sd1)))))));
  localparam signed [3:0] p3 = {{(((-4'sd7)|(3'd6))-(3'sd2))},{(4'd1),((4'd4)<(4'd7))}};
  localparam signed [4:0] p4 = (((3'd5)?(2'd3):(-4'sd6))?(!((-4'sd2)?(-5'sd5):(5'sd15))):(!(-(4'd9))));
  localparam signed [5:0] p5 = (({(5'd6),(-5'sd14),(2'sd1)}<<<{(3'sd1),(2'sd1),(4'd7)})&&({(5'd4),(4'd10)}=={(3'd6),(3'd4)}));
  localparam [3:0] p6 = (((2'sd0)<(-2'sd1))>>((2'd2)-(-5'sd8)));
  localparam [4:0] p7 = (|((&(~&(~((4'd4)<=(-2'sd0)))))+(4'd8)));
  localparam [5:0] p8 = (|(+(|(5'd16))));
  localparam signed [3:0] p9 = ({1{(((-2'sd0)?(5'd27):(5'sd15))^{4{(5'd1)}})}}==(3'd7));
  localparam signed [4:0] p10 = (~^(-4'sd5));
  localparam signed [5:0] p11 = ({2{{2{(5'd18)}}}}<=(~|{1{(((5'd16)|(-5'sd0))>{2{(5'sd11)}})}}));
  localparam [3:0] p12 = (((2'd1)<(2'd2))>=((3'sd1)>>(-5'sd5)));
  localparam [4:0] p13 = ({4{(3'd4)}}===({(5'd26),(2'sd0)}&&((5'sd11)>(5'sd8))));
  localparam [5:0] p14 = ((&(2'sd0))==(4'd2 * (2'd2)));
  localparam signed [3:0] p15 = (~(|(3'd4)));
  localparam signed [4:0] p16 = (|(|(^((-4'sd5)+(((4'sd3)>(-5'sd3))==(+((4'sd2)>>(5'd1))))))));
  localparam signed [5:0] p17 = ((-3'sd1)>(5'sd10));

  assign y0 = ({3{{(b1&a0)}}}<<$unsigned((-2'sd0)));
  assign y1 = (5'sd12);
  assign y2 = ({1{({4{a0}}==(p9+p13))}}?({3{p17}}?{p12,a2}:{3{a3}}):{4{p14}});
  assign y3 = {4{(b4&a5)}};
  assign y4 = ($unsigned(((a0?b0:b2)===((b5+b3)|(4'd2 * a1))))==(($unsigned(p10)!=(p13?p14:p17))&&((p0^~p12)*(p16!=p13))));
  assign y5 = {1{{3{{$signed(p6),(p3),{a2,p16}}}}}};
  assign y6 = ((6'd2 * (a1!=b2))!==(&(&$signed(a2))));
  assign y7 = ((5'sd11)=={3{p14}});
  assign y8 = (((~&b5)-{1{b3}})^~({4{p17}}&(&b0)));
  assign y9 = {3{(4'd0)}};
  assign y10 = (4'd2 * {p14,p12,b0});
  assign y11 = (~&{(p5?p7:a4),{(b5?p8:a4),{p15,p16,a5}},((a0?a2:b5)===(a3|a3))});
  assign y12 = ((^p3)|(~|p9));
  assign y13 = (&(^((~^(~a1))<<(~&(b5!==b1)))));
  assign y14 = ((~&(|((b4?b5:b1)>>(3'd5))))!=={(a0<b4),(b1?a0:b2),(b1<<a4)});
  assign y15 = ({(a3!==b3)}>>((!a5)>>>(p13>>p10)));
  assign y16 = (-4'sd7);
  assign y17 = ($unsigned((|(b3?b0:p5))));
endmodule
