module expression_00104(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~&(-(~(2'sd1))))<<({(5'd19)}<=(^(5'sd5))));
  localparam [4:0] p1 = ((5'sd15)?((-4'sd7)?(3'sd3):(3'sd3)):{(3'sd1),(5'd14)});
  localparam [5:0] p2 = ((3'd7)>>>(2'sd1));
  localparam signed [3:0] p3 = (&(4'd9));
  localparam signed [4:0] p4 = ((((2'sd1)/(2'd3))|((4'd1)/(3'd2)))?(((5'sd12)?(2'sd0):(2'd1))===((-3'sd2)===(5'sd15))):(((4'sd3)?(5'sd2):(-2'sd0))?((-2'sd1)?(3'd3):(4'd9)):((4'd14)<<<(5'd7))));
  localparam signed [5:0] p5 = ({((3'd4)?(4'sd6):(-4'sd3))}>((5'sd8)?(3'd3):(4'd8)));
  localparam [3:0] p6 = (2'd0);
  localparam [4:0] p7 = {(~((3'sd1)<<(2'd3)))};
  localparam [5:0] p8 = (+{1{(&(^{2{(+{{(4'd12),(-3'sd2),(-5'sd0)}})}}))}});
  localparam signed [3:0] p9 = (5'd14);
  localparam signed [4:0] p10 = {{(~^((5'd28)?(5'sd13):(3'sd1)))},(^{(-2'sd1),(-2'sd1),(-3'sd2)})};
  localparam signed [5:0] p11 = ((&((4'd13)&&(4'd8)))-(+(~(-5'sd14))));
  localparam [3:0] p12 = ({2{{1{(~^(3'sd0))}}}}^~(+{{(5'sd3),(2'sd0),(-2'sd0)}}));
  localparam [4:0] p13 = (((4'sd6)?(2'd2):(2'sd1))?((-4'sd0)<=(2'sd0)):(&(2'sd1)));
  localparam [5:0] p14 = (((2'd3)?(5'd19):(2'd3))?((5'd0)?(-5'sd13):(5'sd9)):{(5'sd9),(5'd13),(2'd3)});
  localparam signed [3:0] p15 = (~|{{(3'sd0)},(~(2'sd0)),((4'sd1)?(3'd4):(-2'sd1))});
  localparam signed [4:0] p16 = (^(|{4{(~|(+(2'd2)))}}));
  localparam signed [5:0] p17 = (((4'd9)<(2'd3))==((4'd1)^(-4'sd0)));

  assign y0 = (4'd5);
  assign y1 = (a0===b5);
  assign y2 = $signed((5'd4));
  assign y3 = (~^{p5,p10,p3});
  assign y4 = (4'd7);
  assign y5 = (-({4{(p17==p6)}}|({(b5===a4)}<={(+(~|p8))})));
  assign y6 = ((b3?a5:a1)!==(^(5'sd14)));
  assign y7 = (~&b3);
  assign y8 = $signed(($unsigned({4{p8}})?(5'd2 * (b0>>p1)):$unsigned((p11?p7:b5))));
  assign y9 = (4'd2 * $unsigned((b0===a4)));
  assign y10 = {p15,a3,a2};
  assign y11 = (p7?a4:b3);
  assign y12 = {((b2<<b1)?$signed((p0>>b1)):({a5,p15}))};
  assign y13 = ((({(|a3)}>={b5,a4})<$unsigned(($signed(b5)!={a5}))));
  assign y14 = {(b5?b5:p0),(p1<=b5),(-{b4,b0,b5})};
  assign y15 = {3{(a3>>>b0)}};
  assign y16 = ((~(4'sd4))?(|(~((3'd5)?{4{p11}}:(5'sd13)))):({3{b4}}?(p12^~p13):(~|b3)));
  assign y17 = ($unsigned({3{{$signed(p0),{3{p16}}}}}));
endmodule
