module expression_00401(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{1{{{(4'd0),(-2'sd0),(3'd4)}}}}}};
  localparam [4:0] p1 = {4{((2'sd1)||(5'sd14))}};
  localparam [5:0] p2 = (5'd31);
  localparam signed [3:0] p3 = {(3'd2),(5'sd10)};
  localparam signed [4:0] p4 = (+{{((2'd2)^~(5'd11))},((-3'sd0)?(3'sd3):(2'd1)),{((4'sd2)<(-4'sd0))}});
  localparam signed [5:0] p5 = {3{((~(2'd2))&&((3'd3)<<<(5'd23)))}};
  localparam [3:0] p6 = (~|(((~|(-4'sd7))?{1{(3'd0)}}:((4'd8)&&(4'd10)))?(((-2'sd1)<=(-3'sd0))+((-5'sd11)==(4'd11))):(&{3{(-4'sd0)}})));
  localparam [4:0] p7 = {((3'd7)!==(2'sd1)),(5'd16),{(5'd26),(3'd1)}};
  localparam [5:0] p8 = ((+(&((-2'sd1)<=(-3'sd3))))>(~|(~(~|(&(-5'sd12))))));
  localparam signed [3:0] p9 = {{(4'd13)},((-3'sd2)?(5'sd7):(2'd2)),{(4'sd3)}};
  localparam signed [4:0] p10 = ({1{(3'sd2)}}?{4{(2'sd0)}}:((4'd5)===(3'sd2)));
  localparam signed [5:0] p11 = {4{((4'd3)&&(5'sd2))}};
  localparam [3:0] p12 = (+(4'sd0));
  localparam [4:0] p13 = {(((-3'sd1)<(4'd5))?((3'd7)!==(5'd28)):(5'd1))};
  localparam [5:0] p14 = (3'sd0);
  localparam signed [3:0] p15 = ((3'd1)==={1{(4'sd4)}});
  localparam signed [4:0] p16 = (6'd2 * ((2'd3)>(5'd16)));
  localparam signed [5:0] p17 = (~&((((-4'sd4)?(3'sd2):(5'd3))<(&(2'sd1)))?((-(2'd2))?(~|(5'd12)):((2'd2)>(4'sd4))):((-(-3'sd2))?(|(-4'sd1)):((2'd2)<(-2'sd0)))));

  assign y0 = (^(4'sd4));
  assign y1 = ({p1,a4}?{4{a5}}:{1{{p17}}});
  assign y2 = ((p11>p6)<={p4,p14});
  assign y3 = ((b2-p2)?(p10^~p9):(p8!=p6));
  assign y4 = ({$unsigned(a0),{p13}}?((p5|a2)?$signed(b4):(a2)):{$signed(((+p1)))});
  assign y5 = (p9);
  assign y6 = {1{(~|(-3'sd1))}};
  assign y7 = (~{2{(!(+(|{2{b2}})))}});
  assign y8 = ((a5^~p13)*(b2|p14));
  assign y9 = ((-4'sd2)>>(-(2'sd1)));
  assign y10 = ((5'sd6)>>>((p6?a1:a5)==(a0?b3:a1)));
  assign y11 = (|((!(~&((b2?p9:b3)&(|a5))))<((a4?a5:p7)?(a2!==b2):(a2?a1:a4))));
  assign y12 = (((~p12)%p4)||(~&(~&(~p11))));
  assign y13 = ((!p11)?(a4?a3:p16):(!p8));
  assign y14 = ((-2'sd1)?(p10?p5:p13):(6'd2 * p1));
  assign y15 = (!{(|(|(+(b3<a0)))),(6'd2 * (~&{p13}))});
  assign y16 = ((~^(((+b2)===(!b3))!==((b3<<b3)-(b5||a3)))));
  assign y17 = $unsigned({1{$unsigned($unsigned((-(~&(((p11|b5)|{1{(-p16)}})>((&$unsigned(b5))>>(~^(p10<b2))))))))}});
endmodule
