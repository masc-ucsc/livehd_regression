module expression_00419(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(((+(4'sd0))>={(4'sd1),(5'd26)})?(6'd2 * (~&(4'd1))):{((4'sd2)||(2'sd0)),(~^(3'sd1))}));
  localparam [4:0] p1 = (2'd1);
  localparam [5:0] p2 = {{(4'd2),((3'd3)?(2'd0):(4'sd0)),(2'd1)},(3'sd2)};
  localparam signed [3:0] p3 = ({(&(~^(-3'sd2))),((5'd10)>=(4'd5))}<(&(((4'd14)&&(4'sd3))|{2{(-2'sd0)}})));
  localparam signed [4:0] p4 = (4'd14);
  localparam signed [5:0] p5 = (4'sd6);
  localparam [3:0] p6 = ((((5'd13)|(4'sd2))?((4'd14)&&(3'd4)):((4'd0)<<<(3'd1)))>=({(4'd8)}>(-3'sd2)));
  localparam [4:0] p7 = ((((2'sd0)-(2'd2))?(3'd3):{3{(2'd3)}})&&(2'd3));
  localparam [5:0] p8 = (~^(&(((-(~(-3'sd0)))||(&((-5'sd12)!=(4'd0))))<=(((-3'sd0)!==(2'sd1))===(-(~&(3'sd2)))))));
  localparam signed [3:0] p9 = (((-2'sd0)||(4'd8))^~(~|(5'd9)));
  localparam signed [4:0] p10 = (((-4'sd6)<<<(4'd3))^((5'd27)>>>(3'sd1)));
  localparam signed [5:0] p11 = (-(~&{(2'd0)}));
  localparam [3:0] p12 = (3'd1);
  localparam [4:0] p13 = {4{(5'd4)}};
  localparam [5:0] p14 = (((4'd8)?(5'sd4):(3'sd0))?((2'd3)?(5'd5):(-2'sd0)):((-3'sd2)&&(5'd0)));
  localparam signed [3:0] p15 = {((-3'sd1)?(3'sd2):(2'd0)),{(-4'sd5),(5'd4),(4'sd6)}};
  localparam signed [4:0] p16 = (^(+(~((^(-2'sd1))>(~(-3'sd0))))));
  localparam signed [5:0] p17 = (-5'sd14);

  assign y0 = ((-4'sd5)&(((2'd2)!=(~|p11))==(~|(~|(a2!==a2)))));
  assign y1 = (p13?p17:p1);
  assign y2 = (~&(~|{3{((a5>=b1)?(b2>>>p10):{4{b3}})}}));
  assign y3 = (-4'sd3);
  assign y4 = $signed((~|$signed($signed((+(~^((+(^(~|(+$unsigned((|(!(-p8)))))))))))))));
  assign y5 = ({(&b1),{b2}}-(+(a0&&b4)));
  assign y6 = (3'd6);
  assign y7 = (+(|(|{b4,b2})));
  assign y8 = ($signed((((p0>=p9)|$signed(a4))|$unsigned((b0!=p7))))&&({(b3<<<a4),$signed(a3)}<=($unsigned($unsigned({p17})))));
  assign y9 = ((^(((p13>=p13)<=(p5&p14))^~((+b4)|(p8<p1))))<<<(!{((a0<<a4)==(b5-a4)),$signed((b4==b2))}));
  assign y10 = (2'sd1);
  assign y11 = {(b4==b0),{1{a3}}};
  assign y12 = {(3'sd1),((p5|p6)>>{1{p17}}),{3{p6}}};
  assign y13 = (^{{(b0||p14),(a3!==a0)},{{a0,a3},(p6<<<b5),(b1||a0)}});
  assign y14 = ({2{(4'd13)}});
  assign y15 = {3{{4{a1}}}};
  assign y16 = (~&a3);
  assign y17 = (^(~&{1{(~(~((-(~^{4{a1}}))<({3{p14}}==(b4!=b2)))))}}));
endmodule
