module expression_00952(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((-5'sd4)===((2'd2)|((3'sd2)+(5'd31))))};
  localparam [4:0] p1 = (2'd3);
  localparam [5:0] p2 = ((-5'sd10)>=(((-2'sd0)===(3'd3))*((4'd11)|(5'sd11))));
  localparam signed [3:0] p3 = (((~|(3'd1))?((3'd4)?(3'd4):(-3'sd3)):(~(4'd10)))||((~^((5'sd12)>(-2'sd0)))^((2'd1)?(2'sd0):(4'sd0))));
  localparam signed [4:0] p4 = (4'd2 * ((5'd2)<<<(2'd3)));
  localparam signed [5:0] p5 = {{2{{(4'd10)}}},({(-2'sd0)}>(~&(2'd1))),(((3'sd3)>(4'd4))!={(2'sd1),(5'd24),(-2'sd1)})};
  localparam [3:0] p6 = {4{{1{(-2'sd1)}}}};
  localparam [4:0] p7 = (((5'sd3)?(5'd1):(4'd5))?(4'd13):((-4'sd7)^(-3'sd0)));
  localparam [5:0] p8 = ((((2'd2)?(3'd7):(5'd17))^(&(4'sd5)))!==((3'sd3)?(4'd10):(3'd1)));
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = {(3'd3),(3'd0),(3'sd1)};
  localparam signed [5:0] p11 = ((((3'd5)?(-2'sd1):(-3'sd3))?(4'd6):((3'd2)>=(-2'sd1)))?(((-5'sd9)?(3'sd0):(3'd0))?((3'd5)+(4'd11)):(5'd8)):(((4'd7)^(3'd6))<(5'sd11)));
  localparam [3:0] p12 = {({4{(4'd14)}}<<<{2{(3'd7)}}),(((2'd0)&&(-2'sd1))==((3'd1)^~(4'sd2))),({4{(5'sd15)}}&{(-5'sd3)})};
  localparam [4:0] p13 = ((((2'd1)+(-3'sd2))-((3'sd1)&(5'd17)))&&(((3'd0)-(4'sd7))&&((2'd1)^(-2'sd0))));
  localparam [5:0] p14 = ((3'sd3)?(2'd0):(5'd11));
  localparam signed [3:0] p15 = {4{(-3'sd2)}};
  localparam signed [4:0] p16 = (({4{(5'd9)}}<<<(-(5'sd14)))>>{1{{1{(-(-4'sd0))}}}});
  localparam signed [5:0] p17 = (~|(-3'sd2));

  assign y0 = (~&(^(-$unsigned((((^(a5^~b0))^(^$signed(p10)))&&((~|(a3<<<b1))^(a2>>b3)))))));
  assign y1 = (4'sd5);
  assign y2 = (-3'sd1);
  assign y3 = (2'd0);
  assign y4 = ((-(p11+p6))*(4'sd4));
  assign y5 = (~&((^(~^((~^p13)>{4{p5}})))|((p2>>>p2)?(-p4):(p12&&p9))));
  assign y6 = ($unsigned(({$signed(b0),$signed(p11)})));
  assign y7 = ((|(^((a3>=p12)&(a1+p9))))^((b3<=p16)+(p4*p7)));
  assign y8 = $signed((&((a3?a4:a2)^(b3?b1:a2))));
  assign y9 = {1{{2{(5'd24)}}}};
  assign y10 = (((p5<<p11)/p11)&&(&(&((p16?p14:p15)?(b1?p7:p14):(p6<<<p12)))));
  assign y11 = $unsigned((-3'sd2));
  assign y12 = (3'd7);
  assign y13 = (-(~^($signed(((~(&p17))?{1{{p3,p12,p12}}}:(!(5'd2 * p8))))&({1{((p13>p13)?(p4?b3:b3):(a4<=p6))}}))));
  assign y14 = {{{{b5},{p0}}},{{{b3},{a4,a2}}}};
  assign y15 = (p6?p10:p4);
  assign y16 = ((((a0?b5:a2)&&($signed(b2)<=(b5||b1)))===(^((|(~&(~b3)))-$signed((a2!==a2))))));
  assign y17 = (-(&((b1^~b5))));
endmodule
