module expression_00149(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!{2{(~^(-(~&(~^{4{(3'd5)}}))))}});
  localparam [4:0] p1 = (~((~^((5'd5)^(2'd3)))?((4'd9)?(2'd1):(2'd1)):((-4'sd6)?(4'd7):(3'd6))));
  localparam [5:0] p2 = ((-2'sd0)|(2'd2));
  localparam signed [3:0] p3 = ({2{((-4'sd3)||(4'd9))}}<<<{3{((2'sd0)<=(-3'sd2))}});
  localparam signed [4:0] p4 = (5'sd9);
  localparam signed [5:0] p5 = (((5'sd13)==(3'sd3))?((5'd18)>>>(5'd31)):((4'd11)?(3'd4):(3'd3)));
  localparam [3:0] p6 = {{(-4'sd1),(5'd19),(2'sd0)},(+(!(2'd1))),((4'sd1)<<(-5'sd11))};
  localparam [4:0] p7 = (^((&((5'd9)||(3'sd2)))?({(3'd1),(5'd24)}!={(4'd12),(5'd1)}):((-(4'd1))===((2'sd1)?(-3'sd0):(3'd3)))));
  localparam [5:0] p8 = (((2'sd1)&(3'd4))!=((-2'sd0)?(-3'sd0):(3'd2)));
  localparam signed [3:0] p9 = ((~({1{((5'sd14)>=(2'd3))}}<=(^((-3'sd1)<<<(2'd2)))))&&((((3'd4)>>>(5'd8))||((3'sd2)<<<(2'sd0)))<(&((3'd1)==(4'sd3)))));
  localparam signed [4:0] p10 = (~&(5'd18));
  localparam signed [5:0] p11 = {2{(((4'd11)-(-3'sd2))?((-5'sd2)>>>(3'sd2)):((4'sd2)===(-2'sd0)))}};
  localparam [3:0] p12 = ((^((3'sd3)>(-4'sd0)))<(|(~|{3{(-5'sd14)}})));
  localparam [4:0] p13 = ({2{(((3'sd1)|(5'sd8))>>((2'sd0)>>(5'sd4)))}}>>>({2{((2'sd0)&&(3'd1))}}>(-5'sd0)));
  localparam [5:0] p14 = (3'd2);
  localparam signed [3:0] p15 = (((4'sd6)?(2'sd0):(2'd1))&(-(3'd1)));
  localparam signed [4:0] p16 = (5'd12);
  localparam signed [5:0] p17 = (~|((((5'd2)?(5'sd13):(-2'sd0))===((4'd12)*(3'd7)))+((3'sd0)>=(~(3'sd1)))));

  assign y0 = (5'd6);
  assign y1 = ((~&(~|((b5^~p14)^(b0&&b1))))<<$unsigned((-(|$unsigned((+($unsigned(a5)!==(b2+b2))))))));
  assign y2 = $signed($unsigned(((a0!=p0)<($unsigned(b4)))));
  assign y3 = {(|(~^{4{(&(~&(6'd2 * b2)))}}))};
  assign y4 = (3'd5);
  assign y5 = (((({p13,b3}||$signed(b0))^((p12?p4:p1)<<<$signed(p8))))-(((p16&a4)^~{a4})&&{$signed(b4),{p8}}));
  assign y6 = {1{(((p11&&p3)+(-5'sd7))||{p14,p17,p5})}};
  assign y7 = (-(~^((p10?p2:p7)<<(&p13))));
  assign y8 = ({2{(b3<=b4)}}!==((a5|a1)|{1{(a4<<a1)}}));
  assign y9 = ((-3'sd1)>(((b5>p16)&&(b0>>a0))&&((~b2)+(~&a4))));
  assign y10 = ((+((b3)===(a4>a0)))<<(!(|(a3/p0))));
  assign y11 = (~^(-3'sd1));
  assign y12 = $signed((|(!{2{$signed({(^p15),{p14}})}})));
  assign y13 = (3'd0);
  assign y14 = ((p14>p2)>>{p15,p10,a0});
  assign y15 = (+$unsigned(((((p13<<p6)&(~|p7)))?((4'sd7)?(p15?p1:p10):(p9<=p11)):((b2?p16:p1)?(p13?p2:p2):(|p16)))));
  assign y16 = (&(((!$signed((+((~|p4)<=(5'd14)))))<<<(+((p0<<p2)|(5'sd10))))));
  assign y17 = ((~&p17)>(p5?p3:p13));
endmodule
