module expression_00039(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-(5'd0))&&((2'sd0)?(5'd6):(-2'sd1)))?((3'd5)?(5'sd2):(-2'sd1)):(~^(3'd1)));
  localparam [4:0] p1 = (((-4'sd7)!==(-2'sd0))?((-2'sd1)<<<(2'd2)):((4'sd1)?(3'd7):(-2'sd1)));
  localparam [5:0] p2 = {{(4'sd3),(-5'sd3)}};
  localparam signed [3:0] p3 = (((5'd11)?(3'd3):(-3'sd3))==(5'sd8));
  localparam signed [4:0] p4 = {3{((5'sd0)>=(2'd2))}};
  localparam signed [5:0] p5 = ((-(((2'sd0)>>(-3'sd2))%(-5'sd15)))<(!(((-3'sd3)^(4'd5))>>((5'd10)>(2'sd1)))));
  localparam [3:0] p6 = (~|{(5'sd12)});
  localparam [4:0] p7 = (3'd5);
  localparam [5:0] p8 = {{(4'd5),(-4'sd7),(-5'sd14)}};
  localparam signed [3:0] p9 = (~(+((|(~^(!(^(3'sd3)))))>>>((&(5'd5))||(5'sd2)))));
  localparam signed [4:0] p10 = ((6'd2 * (4'd10))&((2'sd0)!=(3'sd2)));
  localparam signed [5:0] p11 = (2'sd1);
  localparam [3:0] p12 = {2{(5'sd9)}};
  localparam [4:0] p13 = ((&((-5'sd10)<<<(4'd3)))%(-2'sd1));
  localparam [5:0] p14 = ((^{4{(-2'sd0)}})^~(^{3{(2'd0)}}));
  localparam signed [3:0] p15 = (|(3'sd1));
  localparam signed [4:0] p16 = (((-3'sd1)?(4'd13):(-4'sd2))?((3'sd0)?(3'd5):(3'sd1)):((3'sd1)?(-4'sd6):(4'd11)));
  localparam signed [5:0] p17 = (~{(~(~(&{(~|{{3{(-4'sd7)}},(~&{2{(-5'sd0)}})})})))});

  assign y0 = (4'd9);
  assign y1 = {2{((~&a3)==(a2?a0:b1))}};
  assign y2 = (((+(-5'sd4)))>>>$unsigned((-2'sd0)));
  assign y3 = ((~((+(6'd2 * b1))+(-5'sd3)))>>(5'sd5));
  assign y4 = ({({4{a1}}===(b1&a4))}<<{{p12,p17,p2}});
  assign y5 = (!{((a5?p2:p14)>={b4,p9})});
  assign y6 = ((p13?p12:b4)?((p6?b4:b2)<<<(p1?a4:p9)):((p15!=p5)!=(|a5)));
  assign y7 = ((-3'sd3)-((a3?b2:b5)>>>((b4<<<b1)>>(b2^a1))));
  assign y8 = {($unsigned(a4)<={b3,b4,a1}),$unsigned(((&a3)<=(b2>>>p2))),((!b0)>>(~^a3))};
  assign y9 = ((4'd5)-(5'sd6));
  assign y10 = (^{1{((+(|(!(-((~p16)&(+a3))))))<=(~|(((p13!=p9)^(&p14))<<(4'd2 * (~p14)))))}});
  assign y11 = ((3'sd1)?$signed(p7):(a5));
  assign y12 = (((a4?b3:a0)>{a5,b3,b0})!==((5'd2)?(b1|b0):(+a1)));
  assign y13 = $unsigned((-3'sd1));
  assign y14 = (-2'sd1);
  assign y15 = (~{({3{(p3>=b2)}}==(|(~&(!(p5>p8)))))});
  assign y16 = {3{(p3==p5)}};
  assign y17 = (!{a4,b4,a2});
endmodule
