module expression_00805(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(~&(-2'sd0)));
  localparam [4:0] p1 = (!(+(4'd8)));
  localparam [5:0] p2 = {2{(5'd5)}};
  localparam signed [3:0] p3 = {3{(-3'sd2)}};
  localparam signed [4:0] p4 = {{((-5'sd2)?(3'd6):(-3'sd3)),((4'd2)<<(-2'sd0))},{{(5'd2)},{(-3'sd3),(4'd5)},((3'd6)^(4'd11))}};
  localparam signed [5:0] p5 = ({2{(3'sd0)}}+((5'sd1)+(5'sd3)));
  localparam [3:0] p6 = ({1{{((-2'sd1)?(5'd21):(-2'sd1)),((2'd2)^(3'd7))}}}<={{(4'd0),(5'd21),(-4'sd3)},((5'd1)>=(2'd1))});
  localparam [4:0] p7 = (((!(2'd0))&&((-5'sd12)<=(5'd0)))<<(((-4'sd4)>>>(2'd2))^((5'd17)<<<(3'sd2))));
  localparam [5:0] p8 = (((2'd3)>>>(-5'sd8))!=((3'sd0)>(-5'sd2)));
  localparam signed [3:0] p9 = (~((5'd26)-(-2'sd0)));
  localparam signed [4:0] p10 = (!((5'sd7)*(~^((2'd1)?(3'sd3):(3'd6)))));
  localparam signed [5:0] p11 = (&(4'd15));
  localparam [3:0] p12 = {{({2{(2'd2)}}^{(-4'sd5),(-3'sd3)})},{{3{(-4'sd6)}},{{3{(2'd1)}},{2{(5'd27)}}}}};
  localparam [4:0] p13 = (~&((~^({3{(4'd15)}}-{2{(-2'sd1)}}))>={2{((4'd3)<<<(3'd4))}}));
  localparam [5:0] p14 = ((-4'sd2)|(2'd0));
  localparam signed [3:0] p15 = (((4'd12)<<<(2'd1))==((-3'sd3)^(2'sd0)));
  localparam signed [4:0] p16 = ({4{(4'd1)}}!=(^((-2'sd0)^~(-4'sd7))));
  localparam signed [5:0] p17 = {{{3{(2'd1)}},{(-5'sd6),(-2'sd1),(-4'sd1)}}};

  assign y0 = ((5'sd8)<<<(4'd3));
  assign y1 = ((((a1)?(a1==a3):{2{a0}})?{(a5?a0:a5),{b0,a4},{b0,a2}}:({b5,b2}<<{b3,p2})));
  assign y2 = $unsigned(a3);
  assign y3 = (((p5/a0)?(b1<p7):(b5>>>b2))&((b2&p15)<<<(^(5'd2 * p6))));
  assign y4 = (((b0?p8:a4)>>{2{a0}})?({(a1&a3)}>{2{b3}}):((b4?a4:a2)?(4'd14):(a1?p7:p8)));
  assign y5 = ((-$signed((a3?p16:p16)))&&(|(~^(!b2))));
  assign y6 = (((p2<=b5)==(~(~|p3)))+(&(|((a4)%a3))));
  assign y7 = ({2{(b5?b0:a4)}}?((a1?p9:b5)>(~|(a1===b2))):(5'd3));
  assign y8 = $unsigned({{(-(-{a3,b3,a0}))},$signed((~^{p10,p16,p16}))});
  assign y9 = (((~|{4{p15}})!={2{p8}})<((a4>>b5)!==(b1>>>b2)));
  assign y10 = ((p2-b0)+(p3-p13));
  assign y11 = {4{((-p17))}};
  assign y12 = (|$signed((3'd2)));
  assign y13 = ((-(a3*b5))-(~&(b1+a1)));
  assign y14 = (((a1==a1)|(p0<p14))<=((p15!=p1)!=(b2-p6)));
  assign y15 = (({a0,b4,b4}>=(4'd13))?{2{(b2>a0)}}:{{{a3}},(b2?a2:a4)});
  assign y16 = {4{(~(|p2))}};
  assign y17 = (3'd3);
endmodule
