module expression_00482(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd2);
  localparam [4:0] p1 = (+(&(!({1{{4{(2'sd1)}}}}>>>({3{(3'd1)}}>>((3'd3)>>>(5'd16)))))));
  localparam [5:0] p2 = (|(-2'sd0));
  localparam signed [3:0] p3 = ((2'sd1)===(3'd2));
  localparam signed [4:0] p4 = (&(-(3'sd3)));
  localparam signed [5:0] p5 = ((3'sd0)?((-5'sd5)?(2'sd1):(-4'sd7)):(-2'sd0));
  localparam [3:0] p6 = (~^(((-5'sd14)&(4'sd4))+((4'd10)-(-3'sd1))));
  localparam [4:0] p7 = (&(3'd7));
  localparam [5:0] p8 = (~^(((-(3'd4))===(!((3'sd2)==(2'd1))))^~((+(2'd1))>(+(!(2'd3))))));
  localparam signed [3:0] p9 = (~&((~^{(+((2'd1)==(3'd5))),((2'sd0)&(4'sd2))})<<<({((4'sd0)|(2'd3))}^((2'sd0)<=(5'd5)))));
  localparam signed [4:0] p10 = ({(4'd13),(3'sd1),(5'd10)}+(((3'sd2)+(2'sd1))^~((5'sd11)&(-4'sd0))));
  localparam signed [5:0] p11 = {{4{{(4'd11),(3'd0)}}}};
  localparam [3:0] p12 = (4'sd0);
  localparam [4:0] p13 = ((-((4'sd7)?(5'sd9):(3'd2)))?(!{3{(5'd8)}}):(~&{4{(-2'sd1)}}));
  localparam [5:0] p14 = {((((2'sd1)?(2'd1):(2'd0))&((3'sd0)==(-4'sd5)))==={((-5'sd2)&(-2'sd1)),((5'd24)<(4'd15))})};
  localparam signed [3:0] p15 = ({(-5'sd8),(5'sd7),(-2'sd0)}>((4'd2)<(3'd4)));
  localparam signed [4:0] p16 = {2{(-4'sd7)}};
  localparam signed [5:0] p17 = (((-5'sd4)<<(5'd16))^~(3'd0));

  assign y0 = (&p0);
  assign y1 = $unsigned(((a1<p8)&&(4'd2 * a2)));
  assign y2 = {4{{2{a5}}}};
  assign y3 = (+(^(&(~&(~^{4{(|p17)}})))));
  assign y4 = (3'sd0);
  assign y5 = (5'd0);
  assign y6 = (|({3{(~(b0!==a2))}}<={3{(a1||a3)}}));
  assign y7 = (6'd2 * (p2?p14:p1));
  assign y8 = ((^(((a3!==a4)|(b5>p14))!=((+a0)!==(!b1))))>=(((p11>=p3)>>>(p9==p8))<(|(~^(!p16)))));
  assign y9 = (((-4'sd5)>{3{{a2,b3,b5}}})>>(({2{a0}}<=(p4<<b2))!=(3'sd1)));
  assign y10 = (|((p4<<b1)>(p4<<<p1)));
  assign y11 = (p12<<<p4);
  assign y12 = (6'd2 * (b2?b0:b2));
  assign y13 = (({2{(p15?p10:p17)}}<<{1{(b4==a2)}})-{{{(3'sd2),(p1||p15),(!p8)}}});
  assign y14 = (-4'sd0);
  assign y15 = ((p5?b0:b3)<<{(b1?b0:a3),(p4>=a1)});
  assign y16 = (3'd5);
  assign y17 = {(!((+(|(-p0)))<<(3'd5)))};
endmodule
