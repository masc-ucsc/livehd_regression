module expression_00440(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd1)%(-2'sd1))%(-5'sd2));
  localparam [4:0] p1 = {1{{3{(~&((-5'sd5)>>>(4'sd3)))}}}};
  localparam [5:0] p2 = ((^((-3'sd0)>>>(-5'sd8)))||{((-5'sd7)!==(3'd2))});
  localparam signed [3:0] p3 = (~(-2'sd0));
  localparam signed [4:0] p4 = {1{({{(-2'sd0),(-5'sd10),(-5'sd3)}}^(4'd2 * (5'd21)))}};
  localparam signed [5:0] p5 = (&((((4'd14)^(4'd3))^~((-3'sd3)===(3'd1)))^((~(4'sd4))&((5'd10)&(2'sd0)))));
  localparam [3:0] p6 = {(-5'sd4),(2'd2)};
  localparam [4:0] p7 = ({(5'sd8),(2'sd1)}<<(~^(+(2'd2))));
  localparam [5:0] p8 = {(&((~|(4'sd7))&{2{(5'd10)}}))};
  localparam signed [3:0] p9 = (4'sd0);
  localparam signed [4:0] p10 = (3'd2);
  localparam signed [5:0] p11 = {(((5'd7)>>(-3'sd1))||((-3'sd1)&(3'd5)))};
  localparam [3:0] p12 = (|(~&((3'd0)?(2'd2):(3'd3))));
  localparam [4:0] p13 = (!(((3'd5)?(4'd8):(2'd0))?(((2'd1)?(-4'sd7):(-5'sd0))||((5'sd10)?(5'd31):(5'sd15))):((-2'sd0)?(5'd7):(2'd1))));
  localparam [5:0] p14 = {4{{((4'd3)+(-3'sd2))}}};
  localparam signed [3:0] p15 = ((6'd2 * (2'd2))&&{1{{1{(-4'sd3)}}}});
  localparam signed [4:0] p16 = {{((~|(3'd4))^~{(2'sd1)})},(|{((5'd30)<(4'd3)),(^(3'd1))}),(-{(+(4'd15)),(&(2'sd0))})};
  localparam signed [5:0] p17 = ({{(5'd27),(3'sd0),(-5'sd7)}}|{({(4'd13),(-2'sd0)}<<((-5'sd8)<<<(3'd1)))});

  assign y0 = {1{(~|{4{(p9?b1:a1)}})}};
  assign y1 = (2'd1);
  assign y2 = ((((a5!==b5)+{p14,p12,p9})!=(&(~&(b3-b3))))<=((6'd2 * (p13-p0))<<<{1{((b5===b1)>>$signed(p17))}}));
  assign y3 = ((-5'sd1));
  assign y4 = ((-5'sd5)<<(4'd5));
  assign y5 = {1{{3{{{{2{a3}},{a0,b4},{3{p6}}}}}}}};
  assign y6 = $unsigned(($unsigned((~&(~(((~&a1))))))-$unsigned((~&($signed(b5)>>(a2?b0:a3))))));
  assign y7 = {2{(~|((^{1{{4{b3}}}})))}};
  assign y8 = (((p12>=b2)%p0)>>(((p13&p2)|(p13^a2))^~(2'd2)));
  assign y9 = (((-2'sd1)==(-5'sd11))<<<(2'd0));
  assign y10 = (|($signed(b5)));
  assign y11 = {3{{4{(!p15)}}}};
  assign y12 = {($signed(p8)),(p7<<p12)};
  assign y13 = $unsigned((((3'sd2))));
  assign y14 = (5'sd12);
  assign y15 = {1{(((4'd2)||(b4^~b5))>>(((2'd3))|(b2>>a3)))}};
  assign y16 = ((5'd2 * (a2&&b0))?((~(p13<b0))|(p13<=p10)):(!(~&(~|(~&{4{b3}})))));
  assign y17 = {{{{p10,b2,a4},{a4,a3,p7},{{p6,a2,p7}}}}};
endmodule
