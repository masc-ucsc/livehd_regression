module expression_00680(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(-4'sd5)}};
  localparam [4:0] p1 = (6'd2 * ((5'd16)===(4'd6)));
  localparam [5:0] p2 = ((-3'sd3)+(4'sd2));
  localparam signed [3:0] p3 = ((!((4'sd4)+(5'sd11)))||(&((3'd0)&(2'sd0))));
  localparam signed [4:0] p4 = {{(&(!(-(-2'sd1))))},(((3'd5)!=(-3'sd2))^(|(3'd3)))};
  localparam signed [5:0] p5 = ((4'd2)!==(4'sd0));
  localparam [3:0] p6 = (3'd3);
  localparam [4:0] p7 = {({(4'sd1),(5'sd4),(2'd0)}>>((2'sd1)|(-5'sd3))),{{(-2'sd1),(5'sd8),(5'd28)}}};
  localparam [5:0] p8 = (5'sd0);
  localparam signed [3:0] p9 = ((((-5'sd0)||(-4'sd2))&&((2'sd0)?(5'd7):(-2'sd0)))?(((2'sd1)&(5'd4))<((3'd4)*(2'd2))):(((4'd7)<<(4'd6))?((2'sd1)+(4'sd3)):((5'sd5)<=(2'd2))));
  localparam signed [4:0] p10 = (((3'd5)>>>(4'sd2))<((4'sd0)<=(5'sd6)));
  localparam signed [5:0] p11 = (2'd0);
  localparam [3:0] p12 = (+(+((((2'd0)+(3'd7))<=(^(2'd2)))===((~^(2'd3))<<(-(-4'sd3))))));
  localparam [4:0] p13 = {(!((-2'sd1)>>>(3'd1))),(!((4'd15)<<(-2'sd1))),{(5'd28),(2'd1),(-2'sd1)}};
  localparam [5:0] p14 = (((~|(-5'sd14))!==(4'd2 * (4'd15)))<=(((2'd1)?(-2'sd1):(-2'sd0))+((-4'sd4)===(5'sd2))));
  localparam signed [3:0] p15 = ((+(4'd3))?((2'd1)?(5'd17):(2'sd1)):(~^(-5'sd15)));
  localparam signed [4:0] p16 = (~((4'd2)?(~|((-5'sd4)+(2'd0))):(~^(~^(5'sd11)))));
  localparam signed [5:0] p17 = (((4'd8)>>>(2'd2))?((-2'sd0)===(4'd4)):((4'd8)?(3'sd1):(-5'sd3)));

  assign y0 = $signed((($unsigned((|p11))%p16)<<<((b5!==a4)|(b3===b4))));
  assign y1 = (~|p17);
  assign y2 = (~&(!(((p1+p13)&&(~|(-p16)))&&((p12>p4)>>>(!(p12==p12))))));
  assign y3 = (~&(p6?p8:p8));
  assign y4 = (3'd6);
  assign y5 = (~(3'd1));
  assign y6 = (((~|{{1{p0}},{2{p13}}})>>(6'd2 * (&(+p0))))>{(p2+p9),{2{a0}},{(p0?p7:p13)}});
  assign y7 = ((&$signed((&((p11&&p6)^(&p2)))))||(((!b4)^$signed(b0))!==($unsigned(a1)<=(b0<<<b5))));
  assign y8 = {4{(p6||p5)}};
  assign y9 = $unsigned({3{p15}});
  assign y10 = {4{p6}};
  assign y11 = (4'sd5);
  assign y12 = ((-p7)?(-2'sd1):$signed(p7));
  assign y13 = (b2?p2:p5);
  assign y14 = (~|{3{(^(a3^~p13))}});
  assign y15 = ((p15?p5:p1)^(p14>=a4));
  assign y16 = ((a2<<<a1)!=(~&(a5<<a1)));
  assign y17 = {2{$signed((b2>=p0))}};
endmodule
