module expression_00519(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(&((5'd20)?(3'd4):(-2'sd1))),(+(5'sd13)),{(2'd0),(3'sd0),(4'd12)}};
  localparam [4:0] p1 = (4'd6);
  localparam [5:0] p2 = (~^(^(4'd9)));
  localparam signed [3:0] p3 = (~(~&{3{(+(!{3{(5'd19)}}))}}));
  localparam signed [4:0] p4 = (&(~|(((4'd12)?(4'd2):(2'd2))?(~((3'd4)?(-5'sd10):(5'sd10))):((6'd2 * (5'd17))>=((2'sd1)>=(5'd18))))));
  localparam signed [5:0] p5 = ((((4'd2)<<<(3'sd1))==((-2'sd1)&&(2'd3)))>>((5'sd12)<<((3'd6)<=(4'd14))));
  localparam [3:0] p6 = (&(!(((2'd0)!=(5'sd0))?(+(3'd1)):((-2'sd1)<<(2'd0)))));
  localparam [4:0] p7 = ((((2'd1)%(-4'sd7))|((5'd11)^(3'd3)))>>(((-5'sd5)^~(4'sd4))==((-4'sd6)|(2'sd0))));
  localparam [5:0] p8 = {3{(|(3'sd3))}};
  localparam signed [3:0] p9 = {3{(-4'sd2)}};
  localparam signed [4:0] p10 = ((((-4'sd1)?(3'd0):(2'd0))+((-2'sd1)^(3'd2)))<=(((5'd25)!=(4'd14))+((5'sd6)===(-4'sd2))));
  localparam signed [5:0] p11 = (3'd3);
  localparam [3:0] p12 = (!(((4'sd3)-(-5'sd0))===((5'sd15)<=(4'd3))));
  localparam [4:0] p13 = (6'd2 * (5'd17));
  localparam [5:0] p14 = (((-5'sd1)<<<(2'sd1))/(-4'sd0));
  localparam signed [3:0] p15 = ({1{(4'sd0)}}<=((^(4'd1))||((-2'sd0)!=(-4'sd4))));
  localparam signed [4:0] p16 = (^(((2'd3)>>(+(-4'sd6)))&(|{(5'd7),(4'd3),(3'd3)})));
  localparam signed [5:0] p17 = ((-(((-3'sd0)|(5'd26))<(!(!(4'd13)))))|(((-2'sd0)|(5'sd8))|((4'sd5)^(2'd0))));

  assign y0 = {2{{1{(5'sd13)}}}};
  assign y1 = {2{({4{b1}}&&{3{a2}})}};
  assign y2 = ($signed(b5)<{4{p3}});
  assign y3 = {(((~|a2)<<{a0})?(&(-(2'sd1))):{{p13},(!a5)})};
  assign y4 = ((&{4{{p8,p3}}})&&(&({p6,p8,p6}>{p7,p12})));
  assign y5 = {$signed({{(b2^p14),(a0<=p4),{p14,p9,p7}},({p17,p6,b2}&(b0>>a5))})};
  assign y6 = ((-(|(4'sd4)))>=(~|((p14<=b1)?(~|p3):(b1>>>p5))));
  assign y7 = (~(+((a5?p6:p17)?(p4?p16:p12):(-(|p5)))));
  assign y8 = {{(b3?b3:b0),(3'd3),(5'd16)}};
  assign y9 = (({a2,p6,p7}<=(p6<p0))>={(5'd18),(6'd2 * p7)});
  assign y10 = (-((5'd2 * (^$unsigned(b4)))===((b4&&b5)?(a3-b3):(b3?a1:b3))));
  assign y11 = (4'd6);
  assign y12 = (|(((p4?p12:a1))?(p11?a2:p10):(p10?p15:p3)));
  assign y13 = $signed(((+(~&((b2!==b1)^(b1!=b1))))-(&(^(|(+$unsigned((p5?p8:b3))))))));
  assign y14 = (({a1,a0}>=(~^p15))=={(+(5'd0))});
  assign y15 = (((a0===a2)?(a2?a1:a5):(a0?a2:b0))^~(({1{p2}}==(p13>>a3))+{2{(p14^b2)}}));
  assign y16 = {4{(5'sd10)}};
  assign y17 = ((((b1?b3:a0)<<(a4==b1))===({3{b4}}+{1{b5}}))>>{2{((b3&b0)>=(b4||b2))}});
endmodule
