module expression_00832(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd1)?(3'd6):(4'sd2))!==((3'd5)>(-2'sd1)));
  localparam [4:0] p1 = ((-4'sd2)>(-5'sd12));
  localparam [5:0] p2 = ((((5'd5)<(4'd9))|((2'd3)?(-4'sd2):(3'd0)))?(((4'sd4)<<<(3'sd3))!==((5'd9)?(4'd14):(5'd9))):(((2'd0)?(3'sd0):(-3'sd3))?((5'd23)|(5'sd15)):((2'sd0)<<<(-2'sd1))));
  localparam signed [3:0] p3 = (((~^{(3'sd0),(-2'sd0)})>>>(|((2'd3)|(4'd1))))+(~|((2'd3)<=(&(3'sd1)))));
  localparam signed [4:0] p4 = (-2'sd1);
  localparam signed [5:0] p5 = (&(((&{(-2'sd1),(4'd8)})<<{(2'd3),(3'd2)})^(((4'd8)>=(2'd0))>>>{(4'd9),(3'd2),(3'sd1)})));
  localparam [3:0] p6 = {2{{2{{2{(4'sd7)}}}}}};
  localparam [4:0] p7 = {((!(2'sd1))^{4{(2'd1)}}),{2{((4'd2)^~(4'sd6))}}};
  localparam [5:0] p8 = ((4'd0)?(-5'sd11):(4'd8));
  localparam signed [3:0] p9 = (3'd6);
  localparam signed [4:0] p10 = {4{(3'sd3)}};
  localparam signed [5:0] p11 = ((4'd11)?(5'd24):(2'd3));
  localparam [3:0] p12 = {((4'sd7)>>(5'sd3)),(!(!(2'd2)))};
  localparam [4:0] p13 = ((|(-{3{(5'd0)}}))!=(+({3{(-5'sd12)}}-(~&(2'sd1)))));
  localparam [5:0] p14 = (((4'sd6)&(2'd3))>(~(4'd12)));
  localparam signed [3:0] p15 = {2{(+(^(~&((5'sd5)-(3'd0)))))}};
  localparam signed [4:0] p16 = ((((4'd4)<(4'sd0))||{3{(3'd2)}})||((~&(2'd1))-{3{(5'd23)}}));
  localparam signed [5:0] p17 = {({(-2'sd0)}?{(-2'sd1),(5'd25),(3'd0)}:{(2'd0),(-3'sd1)}),((5'd18)?(3'd5):((-5'sd0)<<(3'd0)))};

  assign y0 = (((~(-a3))>>>(a4%p1))^~(^((-b4)*(a0?p11:a5))));
  assign y1 = ($unsigned((p16<<<p11))<=(~|(p10^p1)));
  assign y2 = ({3{$unsigned(p3)}}||{3{(p7)}});
  assign y3 = {4{(+(a4-a5))}};
  assign y4 = ((~&((a1!=a0)!=={3{a0}}))+((^(~|a0))>>{2{b2}}));
  assign y5 = {{1{((-4'sd1)|{3{p9}})}},{({4{a2}}==(~(~&p16)))},(!((a2<=b3)^~(^(&b3))))};
  assign y6 = (({b0,a1,a0}!=={$unsigned({b0})})<((&(a5?b0:a4))<=({b0,p0}<<{b0})));
  assign y7 = (~(((6'd2 * b1)/b3)||((p3*a2)>>(a4!==b0))));
  assign y8 = (~(5'd2 * (b1?a2:p8)));
  assign y9 = ((-{(p7?a4:b3),(p5?a4:p16),{p16,a3}})?{{p10},{4{b0}},{2{p6}}}:{{p2,b0},(p16?p9:b3),{p16}});
  assign y10 = (b5||b1);
  assign y11 = (!(+(&(^p11))));
  assign y12 = ((2'd3)^$signed($unsigned(a0)));
  assign y13 = {1{($unsigned((6'd2 * p0))|{1{{4{b5}}}})}};
  assign y14 = {({p13,p1,p10}?(-p12):{p15,p0}),(~&((p17?p6:p11)?(+p13):{p13})),{{p13},{p12,p11},{p12,p12,p0}}};
  assign y15 = (b4>>>b0);
  assign y16 = ((^((a0>=b1)+(p12+p14)))+((a5^a3)===(b5==b0)));
  assign y17 = ((-4'sd2)<=$signed(((p2>=p8))));
endmodule
