module expression_00192(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd2)/(2'sd1));
  localparam [4:0] p1 = (((-4'sd1)===(-3'sd2))===((3'sd3)||(-4'sd7)));
  localparam [5:0] p2 = (4'd12);
  localparam signed [3:0] p3 = {(-2'sd1),(2'd1),{4{(3'sd1)}}};
  localparam signed [4:0] p4 = (((-5'sd4)?(2'd3):(4'd10))?((4'sd7)===(2'd2)):{(-3'sd1),(4'd14)});
  localparam signed [5:0] p5 = (!({((4'sd2)&(3'd0)),((-4'sd4)>(4'd1))}>=({1{(2'd2)}}>{(3'd7),(3'd3)})));
  localparam [3:0] p6 = (-4'sd7);
  localparam [4:0] p7 = (-4'sd4);
  localparam [5:0] p8 = (+{{4{(3'd5)}},({4{(-4'sd0)}}<=(4'd2)),{(5'd29),(5'sd10),(4'd2)}});
  localparam signed [3:0] p9 = {(-2'sd0)};
  localparam signed [4:0] p10 = ((2'd1)<<(4'sd2));
  localparam signed [5:0] p11 = ((-4'sd4)>>>(2'd3));
  localparam [3:0] p12 = {3{(2'sd0)}};
  localparam [4:0] p13 = ((5'd9)?({(2'd1),(-2'sd0)}>={2{(3'd2)}}):((-4'sd1)?(-3'sd2):(3'sd3)));
  localparam [5:0] p14 = {(((2'sd1)!=(-3'sd2))>>{((5'd14)!=(4'd14))}),(((4'sd3)?(-4'sd6):(4'd1))?((2'sd0)?(-4'sd3):(2'sd1)):((2'd2)-(-3'sd2)))};
  localparam signed [3:0] p15 = ((2'sd1)!=(2'd0));
  localparam signed [4:0] p16 = ({3{((3'd7)|(4'd7))}}+(^((|(-2'sd1))>((-4'sd0)?(4'sd1):(-2'sd0)))));
  localparam signed [5:0] p17 = (~^{2{{(-3'sd3),(4'sd7),(-5'sd9)}}});

  assign y0 = ((-2'sd1)?(p4?p15:a2):(3'sd2));
  assign y1 = ((((a5<<<b5)!==(b4<<<b2))-{(3'd0)})>=(-2'sd1));
  assign y2 = {4{(p12<<b1)}};
  assign y3 = (5'sd11);
  assign y4 = (4'sd7);
  assign y5 = $signed((~&(-(-({4{b5}}>(^(|{p1,a4})))))));
  assign y6 = $signed({(p12>p0),(~&p15),(5'sd14)});
  assign y7 = ({((a1?b3:p15)?(p16?p4:p7):{p5,a3})}?(4'sd0):(+(2'd3)));
  assign y8 = $signed((b0&&b3));
  assign y9 = (4'd15);
  assign y10 = ((a4==b2)>>>(5'sd14));
  assign y11 = ($unsigned(((~(~&a5))>=(5'd2 * b2)))!=((a4?b0:b0)?(a4<=b2):(!(a3^~p14))));
  assign y12 = {1{{1{{1{{{2{a4}},(a2>>a0),(a3+a3)}}}}}}};
  assign y13 = $unsigned($signed(((((4'd6)&(5'd3))^$unsigned($unsigned((-3'sd0))))==$signed({3{(-3'sd2)}}))));
  assign y14 = {4{(!a2)}};
  assign y15 = (~^(-(~|a1)));
  assign y16 = ($unsigned(({(p3>>>p16),(p8<<<p13),(p5&p6)}<<<$unsigned($signed({(b1),{p15,p17,p13},(4'd2 * p0)})))));
  assign y17 = {2{$unsigned($signed({b1,a5,p12}))}};
endmodule
