module expression_00052(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((2'd0)>{(3'sd3)})};
  localparam [4:0] p1 = (^(&(~^((!(~^(-5'sd5)))^((5'd0)<<(2'sd0))))));
  localparam [5:0] p2 = (~|((4'sd0)!=(5'sd12)));
  localparam signed [3:0] p3 = ((&((3'd5)-(3'sd1)))<<(~|((5'd6)^~(2'sd0))));
  localparam signed [4:0] p4 = (((3'd7)?(4'd14):(3'd1))!==(((5'd25)>(-3'sd3))!=={(2'd0),(-4'sd6)}));
  localparam signed [5:0] p5 = (((5'd17)*(-2'sd1))/(4'sd4));
  localparam [3:0] p6 = (((5'sd3)^(4'd4))&&(({(-4'sd0)}>>((4'sd1)||(-2'sd0)))===(3'd4)));
  localparam [4:0] p7 = {3{(4'sd5)}};
  localparam [5:0] p8 = (+(2'sd0));
  localparam signed [3:0] p9 = (~&{((3'd3)>>(2'd0)),((5'd1)>>>(-4'sd4)),((-4'sd0)|(2'd0))});
  localparam signed [4:0] p10 = {1{(-4'sd4)}};
  localparam signed [5:0] p11 = (((5'd11)?(-4'sd0):(-2'sd1))||{(2'd3)});
  localparam [3:0] p12 = {2{{((3'sd3)|(5'sd5)),(+(2'd2)),{(4'd14)}}}};
  localparam [4:0] p13 = ({((2'sd1)?(3'd5):(5'sd9))}&{(-3'sd1),(3'd4),(4'd14)});
  localparam [5:0] p14 = {3{{2{(!(-2'sd1))}}}};
  localparam signed [3:0] p15 = ({(2'd0),(5'd4)}|{(-5'sd13),(-2'sd1)});
  localparam signed [4:0] p16 = (~^(|{1{(!(-2'sd0))}}));
  localparam signed [5:0] p17 = (-2'sd0);

  assign y0 = (+{3{(~^(&(3'sd0)))}});
  assign y1 = (~&$signed((2'd1)));
  assign y2 = ({4{(a0)}}>>>((b0>>>a2)-{1{(a1!==a4)}}));
  assign y3 = ((&(~((~(~|p6))<<(p15!=p7))))<<(|((p6==p9)&(~^(p10!=p7)))));
  assign y4 = {{{p4,b0},{p6}},{(-(^b1))},((p7==p16)!=(p12!=b3))};
  assign y5 = ((4'd2 * (b0?b0:b2))?((p2<<b2)?(b5^~p6):(b0?b2:b0)):((p4>>b5)?(a4?p9:a1):(b3?b2:a2)));
  assign y6 = ($signed((-4'sd0))-(+(+(5'sd7))));
  assign y7 = ((((b3))&{2{b5}})>{2{(p1<=b4)}});
  assign y8 = (~&(2'sd1));
  assign y9 = (~^(4'd11));
  assign y10 = (((a4!=a2)===(b4==b3))||({p15}>>{b4}));
  assign y11 = ((~^(p9<=a2))*(!(b1?a4:b1)));
  assign y12 = (!(+({{a3,b0,a1},(a3?a2:b3)}||{{a4,a5,a3}})));
  assign y13 = ((((a0<<a3)^(b1<<<a3))===((b3<a1)^~(a4>>a2)))+(((b5^~b0)!==(a2>>>b4))===((b4&b3)!==(b2^~b5))));
  assign y14 = (({3{a1}}?{2{a4}}:(a5?p7:p5))?{2{{2{p4}}}}:{2{{a2,p0}}});
  assign y15 = {{4{p10}},{b4,a1,p8},(&p1)};
  assign y16 = (&(~^((p8?p12:p7)>>(!(+b4)))));
  assign y17 = ((3'sd3)!=$unsigned((p15>=p8)));
endmodule
