module expression_00177(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd0);
  localparam [4:0] p1 = (~&(+(+(!(5'd12)))));
  localparam [5:0] p2 = {2{((-4'sd7)?(-5'sd5):(5'd24))}};
  localparam signed [3:0] p3 = ((((3'sd1)<=(3'd2))>>((2'd2)>=(2'sd0)))||(((4'd8)&&(2'sd1))&(~^(5'd12))));
  localparam signed [4:0] p4 = ((~&((4'sd7)<<<(-2'sd1)))?(((3'sd0)|(3'd0))<<<{4{(5'sd5)}}):({2{(-5'sd4)}}+((-2'sd1)+(4'd1))));
  localparam signed [5:0] p5 = (-(5'd23));
  localparam [3:0] p6 = (((5'sd12)?(5'd15):(-3'sd1))!==((3'sd0)?(-2'sd1):(5'd25)));
  localparam [4:0] p7 = {1{(^(&(+{4{(5'd27)}})))}};
  localparam [5:0] p8 = (-2'sd0);
  localparam signed [3:0] p9 = (({(-2'sd0),(3'd1),(4'sd7)}|{(4'sd1),(5'd30)})<=(!(~|(~{{(-2'sd0)}}))));
  localparam signed [4:0] p10 = {(-5'sd0),(4'd6)};
  localparam signed [5:0] p11 = ({(3'd2)}?{1{(2'd0)}}:{2{(2'sd0)}});
  localparam [3:0] p12 = ((((3'd7)?(5'sd12):(-4'sd0))?((5'd8)>=(5'd1)):((5'd12)&&(2'd3)))||(((3'd7)<(2'sd0))||{((-5'sd12)>>(5'sd8))}));
  localparam [4:0] p13 = ((((-4'sd4)&(4'd0))?((4'd10)|(-5'sd14)):((2'd0)===(-4'sd4)))&&(((3'd0)>>>(3'd6))?((3'd3)<(5'sd10)):((-4'sd7)>=(-5'sd4))));
  localparam [5:0] p14 = ({(5'd13),(2'd1)}==(5'd2 * (5'd5)));
  localparam signed [3:0] p15 = (((~|((5'd7)>>(4'sd6)))+(5'd9))>={{(4'd13)},{(3'd7),(3'd0)},(&(!(4'd8)))});
  localparam signed [4:0] p16 = (4'sd2);
  localparam signed [5:0] p17 = ({3{(5'd6)}}&&{1{((-5'sd0)<<(-5'sd15))}});

  assign y0 = ((~(((b3<<b2)>=(~|b3))!=={1{(~^(-b5))}})));
  assign y1 = ((2'sd1)>>>(~(2'd3)));
  assign y2 = ({4{p3}}|$signed({1{(p17>p3)}}));
  assign y3 = (^(~^((+(!(~|(b3?b4:a2))))?((a0?p0:a0)?(a3?p3:p16):(~^p15)):(|(-(-(p16?p15:b1)))))));
  assign y4 = (({1{{p15,b1,p11}}}>(!{b5,p15}))<{{1{{1{{2{b5}}}}}},{(&(|p14))}});
  assign y5 = {4{a3}};
  assign y6 = ((5'd10)?(p2?p14:p9):(5'd27));
  assign y7 = {1{{(^p10)}}};
  assign y8 = ((p0?p2:p7)?{2{p12}}:(^p8));
  assign y9 = (-4'sd7);
  assign y10 = {2{(~&({3{p8}}>>>(5'd12)))}};
  assign y11 = (~((!(!(~&$unsigned($signed((~&{2{((4'd2 * b1)>=(|(a2+p11)))}}))))))));
  assign y12 = ({2{(~p1)}}<={2{{a3,p7,p10}}});
  assign y13 = {{p14,p16},{p6,p17}};
  assign y14 = $unsigned((((-4'sd0)>>>$signed((5'd24)))<<(-2'sd1)));
  assign y15 = (!$signed(a4));
  assign y16 = (^(|(((p8?p11:p14)<(p9?a4:p8))==((&(p12<=p3))>(|(+p3))))));
  assign y17 = (((b2>=a0)>>(p10)));
endmodule
