module expression_00348(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{(3'd2)}}>>((5'd2)?(2'sd0):(5'sd5)));
  localparam [4:0] p1 = (((3'd6)?(4'sd5):(4'd2))^~(~|(5'd3)));
  localparam [5:0] p2 = (&((~|(^(!(|((3'd2)^~(5'd8))))))!==(~|(((3'd6)^~(3'd7))>>>(~^(5'd4))))));
  localparam signed [3:0] p3 = ((&(&(-3'sd3)))%(3'd1));
  localparam signed [4:0] p4 = (!{{2{(+{(3'd7),(4'sd5),(2'd0)})}},{1{({(2'd3),(5'd24)}?((2'd1)?(-4'sd6):(5'sd2)):(+(-5'sd15)))}}});
  localparam signed [5:0] p5 = (-2'sd0);
  localparam [3:0] p6 = ({3{{2{(3'sd1)}}}}^~({(2'd2)}<{3{(2'd0)}}));
  localparam [4:0] p7 = {((3'd6)?(2'd0):(2'd0)),((3'd1)?(5'd11):(-2'sd0)),((4'd5)>>>(4'd0))};
  localparam [5:0] p8 = (5'd18);
  localparam signed [3:0] p9 = ((3'd0)<<<(4'd13));
  localparam signed [4:0] p10 = {{(-4'sd6),{{{(5'd18),(4'sd0),(4'sd4)}}}}};
  localparam signed [5:0] p11 = (!(4'sd3));
  localparam [3:0] p12 = {1{(!(3'd5))}};
  localparam [4:0] p13 = ((((5'd6)==(4'd2))&&((5'd10)&&(5'd19)))>>(-4'sd3));
  localparam [5:0] p14 = (|((((2'd2)!=(2'd1))!=(~(4'd1)))|((&(4'd13))+((5'd10)>>(5'd30)))));
  localparam signed [3:0] p15 = {4{((4'd14)^~(4'sd5))}};
  localparam signed [4:0] p16 = (^{(&{{(2'd3)},{(3'd2),(2'd1)}}),{((-4'sd4)===(4'sd2)),(~&(4'sd3))}});
  localparam signed [5:0] p17 = {1{(4'd7)}};

  assign y0 = {(({3{(&b3)}}!=={(a0<=a3),{b1,a2}}))};
  assign y1 = (~((|(p1<<p8))|(|(&(p6*p0)))));
  assign y2 = (|(~^{1{{3{(-{1{(+(p12^~a3))}})}}}}));
  assign y3 = ((((p1&p2)>>>(p3-p6))>>((b2*p17)%p14))!=((a2>p14)?(p2>>p15):(p11?b3:b1)));
  assign y4 = ((p0>>>p7)+(~&p16));
  assign y5 = ((^(&p1))?(|(p7>p14)):(2'd3));
  assign y6 = ({1{{4{a4}}}});
  assign y7 = (-(~&p1));
  assign y8 = ($unsigned(($signed(((a2?b3:b1)?$unsigned(a5):$signed(b0)))?$unsigned(((b3)?(a3):$unsigned(a2))):((a3?a0:a4)?(a2?b0:a1):(b0?b2:a1)))));
  assign y9 = (|(!((p8>=p8)*(p8^~p10))));
  assign y10 = ((p10?b5:p4)?{p0,p12}:(p13?p1:p5));
  assign y11 = {1{{1{((~&$signed({1{(5'd31)}})))}}}};
  assign y12 = ((4'd4)===({(3'd3)}<=({b1,a1}<(3'sd2))));
  assign y13 = ((4'd2 * (b2<=p1))<=($signed(((p8<<<p11)<=(a1>=p1)))|{(b2),$signed(b2)}));
  assign y14 = ((-p16)?(+p8):(!p11));
  assign y15 = (p4?p10:p5);
  assign y16 = {{2{{2{b2}}}}};
  assign y17 = {2{({1{{3{p3}}}}^(6'd2 * (b2!==a1)))}};
endmodule
