module expression_00838(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd6)?(-5'sd14):(2'sd1));
  localparam [4:0] p1 = (|(4'sd0));
  localparam [5:0] p2 = (~((5'sd4)|(-2'sd1)));
  localparam signed [3:0] p3 = (4'd5);
  localparam signed [4:0] p4 = {3{(~&(~^{1{(2'd3)}}))}};
  localparam signed [5:0] p5 = (((-4'sd2)-(4'd13))<<<(^(3'd3)));
  localparam [3:0] p6 = {4{(4'd13)}};
  localparam [4:0] p7 = (^{(((5'd8)<(4'sd4))>>>((3'd5)+(-4'sd2))),(3'd3)});
  localparam [5:0] p8 = (((2'd2)<=(-4'sd3))^((-4'sd5)+(3'd1)));
  localparam signed [3:0] p9 = (-3'sd3);
  localparam signed [4:0] p10 = (3'd2);
  localparam signed [5:0] p11 = ({((4'd11)>(5'd7)),(~&(-4'sd6))}||{3{(-5'sd14)}});
  localparam [3:0] p12 = {(~^{{(3'd5),(-5'sd9),(5'd29)},{((4'sd3)>>(2'sd1))},(~&{2{(-4'sd3)}})})};
  localparam [4:0] p13 = (((~(3'd6))<((-3'sd0)==(5'd4)))^({2{(2'd2)}}==={4{(2'sd1)}}));
  localparam [5:0] p14 = {4{{4{(4'd2)}}}};
  localparam signed [3:0] p15 = ((-5'sd7)>(5'd12));
  localparam signed [4:0] p16 = (~&(+(2'sd1)));
  localparam signed [5:0] p17 = ((3'd0)?(2'd2):((2'd2)<<<((-4'sd6)?(2'd3):(5'sd12))));

  assign y0 = (5'd14);
  assign y1 = (|((p8^~p2)||(p4>>p10)));
  assign y2 = (&{4{(|(|{p9,p9}))}});
  assign y3 = {2{({4{p9}}<<<((p12+p8)==(p15<p5)))}};
  assign y4 = (3'd6);
  assign y5 = (((p15?a1:p0)?(b3?p15:a2):(5'd2 * a0))?((6'd2 * a2)?(p5&b4):(p15!=a4)):((!a1)?(p0<b3):(b5===b4)));
  assign y6 = (a4&&b2);
  assign y7 = (((6'd2 * (b0?b1:a0))&({3{b1}}==(b2>=b1)))!==((6'd2 * (b1>>a2))-(~(+(b0||a0)))));
  assign y8 = ((((~&b4)===(&b5))?$signed({2{p7}}):((p17?b5:a1))));
  assign y9 = ({(!{1{{3{p12}}}}),{$unsigned(((p10<p3)))}}>>>{3{{(p5>=b2)}}});
  assign y10 = ($signed(((-(^($unsigned((p5))==$signed((p12)))))|((p16?p9:p3)>>((~&p11)^(^p15))))));
  assign y11 = ((~&{3{(|p0)}})?{(-(a4?p16:p13)),{{4{a3}}}}:{(-{a3}),{4{b0}}});
  assign y12 = ((^(&{1{(-(4'd2 * p0))}}))||(-4'sd0));
  assign y13 = (p1!=p4);
  assign y14 = (-5'sd7);
  assign y15 = {{p7,p4,p6},$unsigned({$signed(a0)}),{(p10?p1:p17),(4'd0)}};
  assign y16 = ($unsigned(p12)+$signed(p13));
  assign y17 = (((p0>>>a0)^~(p2+p10))?({2{p11}}>>>(p11<a4)):$unsigned((p0<p11)));
endmodule
