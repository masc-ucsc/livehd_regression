module expression_00400(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd4);
  localparam [4:0] p1 = {{3{(2'd1)}}};
  localparam [5:0] p2 = ((((5'd0)*(3'sd0))!=((4'sd5)<<(5'd4)))<=(((3'sd0)^~(5'd2))+((-4'sd3)|(-5'sd9))));
  localparam signed [3:0] p3 = (({(5'd23),(3'sd0)}||{2{(5'sd6)}})^~(~(|((-(-3'sd0))&&{4{(2'sd0)}}))));
  localparam signed [4:0] p4 = ((((3'sd3)===(-5'sd13))==((3'sd2)?(4'sd6):(4'd10)))<<<((~|(4'd3))-(~(2'sd0))));
  localparam signed [5:0] p5 = (~|(&(~&(^{4{(2'sd0)}}))));
  localparam [3:0] p6 = ((^((3'sd0)&&(-2'sd0)))>=((-(2'sd0))>(~(3'sd2))));
  localparam [4:0] p7 = {1{((((-3'sd1)>>(5'd3))?((4'sd3)?(3'd3):(3'sd3)):{1{(2'd2)}})&{3{(+(4'd9))}})}};
  localparam [5:0] p8 = {2{(4'sd4)}};
  localparam signed [3:0] p9 = {4{(~^(5'd2))}};
  localparam signed [4:0] p10 = {(2'd3),{(-3'sd1)},{(-2'sd1),(5'd25)}};
  localparam signed [5:0] p11 = {({4{(-4'sd7)}}?{(-5'sd13),(3'd1),(4'sd4)}:{(2'd0),(3'sd3),(3'd4)}),{((3'sd0)?(-5'sd9):(4'd7))},(((4'd4)|(2'sd0))?{4{(2'sd1)}}:(2'd2))};
  localparam [3:0] p12 = (-((~(2'sd0))?(~(5'd0)):{1{(5'd30)}}));
  localparam [4:0] p13 = (^(~(-4'sd2)));
  localparam [5:0] p14 = (&(((3'd4)<(3'd5))*((-3'sd1)/(5'sd3))));
  localparam signed [3:0] p15 = (((3'sd1)?(2'd1):(5'sd15))?{4{(-4'sd4)}}:((5'sd7)?(4'd1):(-2'sd0)));
  localparam signed [4:0] p16 = ({2{((2'sd0)===(4'sd7))}}+{2{((3'd6)?(-4'sd1):(2'sd0))}});
  localparam signed [5:0] p17 = ((~&(!(~^{3{(2'sd1)}})))>(5'd2 * ((3'd1)^~(4'd0))));

  assign y0 = (!{2{(2'd3)}});
  assign y1 = ((p7||p7)|(|p6));
  assign y2 = {$unsigned((+(a0&&p10))),{(p16?p12:p17)}};
  assign y3 = (|(5'sd6));
  assign y4 = (p4<<a4);
  assign y5 = (!(p12?b5:p10));
  assign y6 = (4'd14);
  assign y7 = ((a1>=b4)?(b4>b3):$unsigned((a5>>b2)));
  assign y8 = ((((a3>p6)|(p14|p13))+{4{p14}})>>>{(({p2,p14}<<<{p3,p14})||((p12<<p16)^{p8}))});
  assign y9 = (5'd2 * {4{p8}});
  assign y10 = (-2'sd1);
  assign y11 = ({{{(b2!==b2)}}}-{{p1,a4,p16},(p8>=b2)});
  assign y12 = (a5>=p17);
  assign y13 = $signed({($signed((p15?b5:p6))?{$signed({4{a2}})}:(p14?p16:a4))});
  assign y14 = {(|((^a5)?(a2):(3'sd1)))};
  assign y15 = ((p3?p14:p10)==(b4>>>p0));
  assign y16 = (6'd2 * {(^p7)});
  assign y17 = (^(($unsigned(p5)?(p7<p10):(p6&&p8))?((3'd0)<{p11,p10}):((p16-p6)?(~|a4):(p14|p9))));
endmodule
