module expression_00066(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{((-5'sd8)<(~^((-3'sd0)>>>(3'sd1))))}};
  localparam [4:0] p1 = ((~((5'sd9)^~(2'd2)))>>{2{(~|(-3'sd1))}});
  localparam [5:0] p2 = {{3{((-2'sd1)?(2'sd1):(2'd3))}},{1{((-2'sd0)?(3'sd2):(3'd4))}},{{(-3'sd2),(-5'sd6)},{1{(5'd17)}}}};
  localparam signed [3:0] p3 = {1{(-(((~|(3'd3))||(-(4'd1)))&(((3'sd0)<<(4'sd0))=={1{(-3'sd2)}})))}};
  localparam signed [4:0] p4 = ((-4'sd2)===(3'd4));
  localparam signed [5:0] p5 = ((2'd1)?(2'd2):(-4'sd7));
  localparam [3:0] p6 = (~&{4{{(3'sd2),(3'd7),(4'sd4)}}});
  localparam [4:0] p7 = {1{{3{((5'sd0)>(2'd0))}}}};
  localparam [5:0] p8 = (&(5'sd12));
  localparam signed [3:0] p9 = ({2{(3'd0)}}+{{2{(4'd9)}}});
  localparam signed [4:0] p10 = (((2'd2)>>>(4'sd0))!={((3'd5)||(3'sd0))});
  localparam signed [5:0] p11 = ({(4'd7),(-5'sd14)}!==((-3'sd2)>(5'sd9)));
  localparam [3:0] p12 = ((-2'sd0)<<{{4{(2'sd0)}}});
  localparam [4:0] p13 = (|(5'sd9));
  localparam [5:0] p14 = {1{(2'd0)}};
  localparam signed [3:0] p15 = (6'd2 * ((2'd1)===(4'd3)));
  localparam signed [4:0] p16 = ((((-3'sd1)>>>(5'sd0))/(2'd0))-(4'd2 * ((3'd3)^(3'd0))));
  localparam signed [5:0] p17 = ((4'd9)||(5'd24));

  assign y0 = {{((-{p15,a2})<<<{a5,a0}),({{3{a2}}}>>($signed(p7))),(((((a3+b0)>>>{a2,a1,b3}))))}};
  assign y1 = ((((4'd2 * p7)>(p4>>p9))>=(({p3}<={2{p15}})))<<<$unsigned($signed((((p13||p7))?(a1>>>p13):{3{p14}}))));
  assign y2 = ($signed((|(~|$signed((&($signed(p10)<=(p4>p4)))))))<<<({$unsigned({a1,a2})}!==({2{a0}}==(~^b5))));
  assign y3 = ((~(!(5'sd2)))<={3{(a3^a5)}});
  assign y4 = (2'd0);
  assign y5 = ((((a1+a2)>>(5'd2 * a1))+({b1}<<<{b4,a1,a4}))!=={({a2}>=(b0!=a5)),{((b3>>b2)+(b2||b4))}});
  assign y6 = (((p7<=p5)*(|p15))?((p9?p6:b3)?(p0>>p11):(-p11)):(2'd3));
  assign y7 = (a5>>b4);
  assign y8 = (b0|p3);
  assign y9 = (((~^(^(~^a3)))+((~a3)>{a1,b1}))>(~^(+{{(!(&{a5,a3}))}})));
  assign y10 = $unsigned((b4&&a2));
  assign y11 = {(4'd2)};
  assign y12 = {$unsigned((({(p14?b0:b5)})?($unsigned($unsigned($unsigned(b0)))):{(b5?a0:p4)}))};
  assign y13 = (~&(((b2===a0)<<<(p0>>>p15))<=((a3==p7)&(p8&&a5))));
  assign y14 = (~|(+a4));
  assign y15 = {2{(~^(-2'sd0))}};
  assign y16 = (!{{1{(p17?a2:p8)}},{2{(b0?a0:b1)}}});
  assign y17 = {(({3{a0}})),$signed(({3{a4}}))};
endmodule
