module expression_00795(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(((-2'sd0)==(5'd27))||((5'sd3)^(-4'sd6)))}-{{(4'd9),(3'd5)},((5'd30)|(5'd17)),((3'sd0)&(-3'sd2))});
  localparam [4:0] p1 = (^(~|(^{{3{(~|(-4'sd2))}}})));
  localparam [5:0] p2 = (-(|{(5'd27)}));
  localparam signed [3:0] p3 = (-4'sd2);
  localparam signed [4:0] p4 = ((((5'd22)>=(2'sd0))===((-3'sd2)>(3'd7)))+(((5'd15)+(-4'sd7))===((-5'sd13)!==(3'sd1))));
  localparam signed [5:0] p5 = (-(((4'd10)?(3'sd1):(4'd6))?{1{((2'd0)^(3'd6))}}:((4'd13)?(5'd12):(5'd1))));
  localparam [3:0] p6 = {(~&(5'sd4)),(3'd7),((4'sd2)^(3'd7))};
  localparam [4:0] p7 = (+(|((+(-4'sd5))!=(2'd2))));
  localparam [5:0] p8 = (-(-(+{4{((3'sd0)>=(5'd30))}})));
  localparam signed [3:0] p9 = {3{(-4'sd2)}};
  localparam signed [4:0] p10 = {4{(~(~(3'sd1)))}};
  localparam signed [5:0] p11 = {{((4'd12)|(4'd8))}};
  localparam [3:0] p12 = (~&((((2'd3)|(2'sd1))===((4'd8)+(5'd7)))|((&(4'd2 * (5'd25)))!==((2'd2)>>(-3'sd1)))));
  localparam [4:0] p13 = (3'sd3);
  localparam [5:0] p14 = ((-4'sd1)|(|((-5'sd5)?(3'd4):(5'd24))));
  localparam signed [3:0] p15 = ({(&{4{(4'd9)}}),((4'd13)?(3'd5):(-5'sd3))}&{((3'd3)===(2'sd1)),((5'd30)?(-5'sd13):(2'sd1)),(-2'sd0)});
  localparam signed [4:0] p16 = (~|((5'd22)?(-2'sd0):(-2'sd0)));
  localparam signed [5:0] p17 = {{{(4'd8),(2'd3)},(|(+(-4'sd3)))},{(~^(^(~|(^(!(-4'sd5))))))}};

  assign y0 = (|(&(|(&(~^(|(~^b3)))))));
  assign y1 = (^((|{{a5,a2},(b5&&a3),(~|{a0,a1,b2})})===({(b1+b1)}&(~|(b3>=a4)))));
  assign y2 = ((~(b5))/a2);
  assign y3 = {3{($signed(p14)?(5'd5):(|p0))}};
  assign y4 = (!(!((p11?a2:p4)?(~(+a4)):(|(~&b5)))));
  assign y5 = $signed(({3{b2}}^~(3'd1)));
  assign y6 = ((&((b1+p15)?(&a4):(p16>=p14)))+$signed($signed(((b3&a3)|(b1||p5)))));
  assign y7 = (!((a1>b1)>=(b0===a1)));
  assign y8 = ({4{b5}}<<{a1,a0,p16});
  assign y9 = {(((b0|p0)>>(a0!==a3))==$unsigned(((p11&a5)>>>(~&(p8==b1)))))};
  assign y10 = (!((&(4'd2 * p14))||(a5>=p15)));
  assign y11 = $unsigned({{4{(b5)}},(!(^(&{2{(^(~^p17))}})))});
  assign y12 = (~^(p14));
  assign y13 = {4{((a5|p11)>>{4{p5}})}};
  assign y14 = (~^(~&(((^(-p1))/p7)&&(+((~|p0)*(p3^a0))))));
  assign y15 = (~|(5'sd7));
  assign y16 = (~^(-2'sd1));
  assign y17 = (3'd5);
endmodule
