module expression_00844(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-((-2'sd1)?(2'd3):(5'd1)))?{3{(-3'sd2)}}:(-3'sd3));
  localparam [4:0] p1 = {{(3'd7)}};
  localparam [5:0] p2 = {((-4'sd4)!=(-3'sd2))};
  localparam signed [3:0] p3 = (^{(((3'd0)&(4'sd2))&&((-4'sd0)>>>(3'sd1)))});
  localparam signed [4:0] p4 = {(^{1{(2'sd0)}}),((4'sd6)<<<((4'd6)?(4'sd3):(2'd1))),({(3'sd3)}?((4'd4)?(5'sd12):(-5'sd10)):((5'sd12)?(-3'sd2):(2'sd1)))};
  localparam signed [5:0] p5 = ((~^((5'sd7)|(3'd7)))||(2'd0));
  localparam [3:0] p6 = ((((2'd3)<<<(4'sd7))||(+(-2'sd1)))!==((-2'sd0)?(5'd2 * (3'd6)):(-(4'd14))));
  localparam [4:0] p7 = (-4'sd3);
  localparam [5:0] p8 = (((-4'sd3)^(5'd17))<<((-2'sd0)|(-5'sd2)));
  localparam signed [3:0] p9 = ({(3'd0),(3'd3)}<((2'sd0)?(5'd25):(4'sd7)));
  localparam signed [4:0] p10 = ((~|(~&(-(^(5'd14)))))^~(&(~|(4'd2 * (3'd0)))));
  localparam signed [5:0] p11 = ((3'd5)===((5'd17)<=(5'd4)));
  localparam [3:0] p12 = ((((2'sd0)<<<(3'sd2))>=((5'd4)!=(2'sd1)))===(((-4'sd6)==(-5'sd12))<<<((2'sd0)>=(5'd30))));
  localparam [4:0] p13 = (+(~|{(~^(2'd2))}));
  localparam [5:0] p14 = (~(~(|(~|(~^(|(-(-(!(+(~&(-5'sd1))))))))))));
  localparam signed [3:0] p15 = (+((3'd7)?(2'd3):(3'd3)));
  localparam signed [4:0] p16 = ((3'd2)<(-2'sd1));
  localparam signed [5:0] p17 = ((2'd1)?(2'sd1):(5'd3));

  assign y0 = $unsigned((((p9!=p7)%b1)<<<((4'd2 * p14)<(p5<p4))));
  assign y1 = (b0>>>b0);
  assign y2 = {{2{{(3'd0)}}},{2{{p13,b1}}}};
  assign y3 = {1{(((p16!=p9)&(b2===b3))>>>((p7^~p4)?(p13<p5):(p1==p17)))}};
  assign y4 = (~^{$unsigned($unsigned((4'd6))),((!a3)!=(|p15)),{p16,p11,a1}});
  assign y5 = (4'sd4);
  assign y6 = {((a4?p5:a3)&$signed(p4))};
  assign y7 = ((^(($signed((p17))?(3'sd3):(p6?p17:a1))))^~((p13^~p1)?(a3?b4:b1):$signed((b5<<a1))));
  assign y8 = {1{((({3{b4}}===(b2!=b1))|((b5<<a5)+(5'd2 * a2)))!=={1{({3{b3}}^(a2>>a5))}})}};
  assign y9 = (((~$unsigned(b3))*(~|(+b5))));
  assign y10 = (|((4'd2 * (p1>=p8))<=((+(|(p13>>p11)))^~$signed((|(p15||p8))))));
  assign y11 = (^(^(({a1}<={p14,p6})=={(+p17),(^p13)})));
  assign y12 = (((|p6)?(p6?p4:p2):(|p17))<<(+($unsigned($unsigned(b3))|{1{(p14>=a2)}})));
  assign y13 = (p3%p10);
  assign y14 = (4'sd0);
  assign y15 = ((!a1)?(a1):(6'd2 * b2));
  assign y16 = (+((a5!==a0)?(b0&p11):(p14<<<p8)));
  assign y17 = $unsigned(($signed(((3'sd2)^{((p13!=p7)>>>{p4,p9,p8}),(&(5'd8))}))));
endmodule
