module expression_00082(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^(+(|(!{(-3'sd1),(!{{(2'sd0)},(~^(4'd11))})}))));
  localparam [4:0] p1 = ((!(-5'sd7))>>>(((-4'sd5)?(5'd30):(2'sd0))<<<((-2'sd1)/(-5'sd10))));
  localparam [5:0] p2 = {3{((~|(2'd0))?(2'd1):(^(-2'sd0)))}};
  localparam signed [3:0] p3 = ((2'd1)?(5'd4):(-2'sd0));
  localparam signed [4:0] p4 = {2{{2{(4'd2 * (3'd7))}}}};
  localparam signed [5:0] p5 = ({4{{(2'sd1),(4'd15)}}}||{((2'd3)>=(3'd1)),((-3'sd0)&(4'd12)),((2'sd0)<=(4'sd2))});
  localparam [3:0] p6 = ((~((^(-2'sd1))/(-5'sd3)))<<<(((-5'sd8)>=(5'sd15))+(5'd0)));
  localparam [4:0] p7 = {4{(-2'sd1)}};
  localparam [5:0] p8 = (((2'd2)?(2'd0):(5'sd11))^{(2'sd1),(2'sd0),(-5'sd6)});
  localparam signed [3:0] p9 = (+(3'd2));
  localparam signed [4:0] p10 = (~&(~^((5'sd6)?(2'sd0):(2'sd0))));
  localparam signed [5:0] p11 = ((2'sd1)?{(2'sd1)}:((-2'sd1)?(-3'sd2):(3'd2)));
  localparam [3:0] p12 = (5'd2);
  localparam [4:0] p13 = ((((5'sd4)!=(2'd3))&&(5'd18))<<<{{(4'd3)},((5'd8)&(4'd13)),(-4'sd3)});
  localparam [5:0] p14 = (+((!(+(-3'sd3)))<=(-5'sd4)));
  localparam signed [3:0] p15 = (~|((&(-4'sd0))&&{(2'd2),(-2'sd1)}));
  localparam signed [4:0] p16 = ((3'd5)<<(5'd17));
  localparam signed [5:0] p17 = (({3{(4'sd1)}}==(((-5'sd11)>(4'd8))^((-4'sd6)+(-2'sd0))))<={1{(((5'sd14)>>(-4'sd4))&{2{(2'd3)}})}});

  assign y0 = ({1{(5'd2 * (p1&p1))}}-{4{(b5?p13:p14)}});
  assign y1 = (3'd1);
  assign y2 = (4'd0);
  assign y3 = ({1{(4'd11)}}<$unsigned((4'd2 * (5'd3))));
  assign y4 = (p1<p3);
  assign y5 = ((~|(p5?p4:b5))?(~(&p3)):(|(&p13)));
  assign y6 = $signed($unsigned((p9)));
  assign y7 = (($unsigned(p0)?(p10<=b1):(~|b1))?{3{{3{p10}}}}:(((p12<=p10))-(6'd2 * p0)));
  assign y8 = $signed((|$unsigned((2'd1))));
  assign y9 = (((a2===b1)>>(p0|p6))?((b5?b1:b3)===(b2!=b2)):((b4&&b0)-(p10!=b4)));
  assign y10 = {$unsigned(($signed({(a3|b4),({p5}),(p10&&b2)})>>$unsigned({(^(+(-b4))),($unsigned({b5,a1,a0}))})))};
  assign y11 = ((((-a5)<(b5>>b1))+(4'd12))!=(~|{4{(b2+b3)}}));
  assign y12 = (2'd2);
  assign y13 = (((~|{1{{4{p15}}}})?(~^(+{p6,p15,b0})):(p0?b1:a1)));
  assign y14 = (~|(((!(~a4))==={4{b5}})^(^((b1<<<a3)-$signed(a3)))));
  assign y15 = (~$unsigned($unsigned($unsigned(((|(p3?b3:b3))?(~&(a3?b4:b3)):(|(b2?b2:b5)))))));
  assign y16 = {{2{($unsigned(p4))}}};
  assign y17 = (~|(+(a3<<p2)));
endmodule
