module expression_00307(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(~(4'd13)));
  localparam [4:0] p1 = ({(5'd18)}===((-5'sd11)<<(3'd2)));
  localparam [5:0] p2 = (((-5'sd9)?(4'd12):(2'd3))>>((4'sd1)^~(-5'sd11)));
  localparam signed [3:0] p3 = (((~((2'sd1)<(2'd0)))>((2'd0)&(5'd27)))+(((-4'sd6)<(3'd0))>=((2'sd1)>(3'sd1))));
  localparam signed [4:0] p4 = (~|(~&(|(4'd2))));
  localparam signed [5:0] p5 = (({3{(5'd1)}}<<<((2'd2)^(5'd30)))=={1{{3{(4'd9)}}}});
  localparam [3:0] p6 = ({2{(5'd20)}}>>>((2'd0)>(2'd2)));
  localparam [4:0] p7 = {{1{((-2'sd1)?(5'sd14):(4'd10))}},((3'd0)?(4'sd5):(3'sd2)),((5'd4)?(5'd20):(-4'sd7))};
  localparam [5:0] p8 = {(5'd0),(4'sd4)};
  localparam signed [3:0] p9 = {2{(|(^(2'd1)))}};
  localparam signed [4:0] p10 = (~^(~(5'd2)));
  localparam signed [5:0] p11 = (((3'd1)?(5'd25):(5'sd12))?((5'd8)?(5'd20):(3'sd3)):((3'sd2)>>(3'd3)));
  localparam [3:0] p12 = (((-5'sd11)&{(-3'sd3),(-3'sd0)})<<<((5'd29)+(5'd2)));
  localparam [4:0] p13 = (((3'd1)===((3'd6)===(5'd29)))===(5'd4));
  localparam [5:0] p14 = {(!{2{((-((-2'sd1)<<<(3'sd3)))>>>((3'd0)?(3'd6):(2'd2)))}})};
  localparam signed [3:0] p15 = (-4'sd1);
  localparam signed [4:0] p16 = {1{{{1{{1{(3'd3)}}}},{2{(-4'sd0)}},{1{(!(5'sd4))}}}}};
  localparam signed [5:0] p17 = (3'd4);

  assign y0 = {(~^(&a0)),(a5<<b5)};
  assign y1 = {2{(((b0!==b5)>(p5>>p4)))}};
  assign y2 = (&{{{4{a3}}},((~|b1)|{4{b0}}),$signed((a5==a4))});
  assign y3 = {(b3?a4:a0),{a0,b4,a5},(a5?a0:a1)};
  assign y4 = (((b3<=p17)-(p10?p4:a2))?((p2<<<p7)/p12):((a1?p11:b0)<<<(p9&a4)));
  assign y5 = (~(~|(&(&(|(&(^(!($signed(((-(!b5)))))))))))));
  assign y6 = (+{2{$unsigned(a4)}});
  assign y7 = (4'd11);
  assign y8 = ((((-3'sd0)||(a2?a5:b5))===(b1?a4:a3))&&((3'sd0)?{1{(5'd11)}}:{{b3,p0,p6}}));
  assign y9 = (&(~|(~{(~|(p14>a5)),(!(&a2))})));
  assign y10 = (-5'sd3);
  assign y11 = (~|{((p11&&p12)>>>{4{a3}}),{4{p14}}});
  assign y12 = $signed({2{p9}});
  assign y13 = $unsigned(((-$unsigned($unsigned((+(p6>>p14)))))?(^{(5'd2 * p0),$signed(a2),(p15?p2:p15)}):$signed((((p12?p16:p13)<<(a3?p8:p2))))));
  assign y14 = (({(a0&&a1)})?(b3?b4:b4):{(b4?p8:a3)});
  assign y15 = ($signed((a3?b0:p7))?((p6>=b3)<<<(p14<<<p6)):((a2?p5:b1)-$unsigned(p11)));
  assign y16 = ((!(+((p11<<a2)>>>(5'd2 * p13))))<(((p2<=b3)<=(p11/a1))!=((p12&&b5)^~(b3^b5))));
  assign y17 = {2{{1{(-4'sd2)}}}};
endmodule
