module expression_00971(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~(!(!(3'sd3))))!==(((4'sd6)>>>(-4'sd2))||((5'd15)?(2'sd0):(5'd30))));
  localparam [4:0] p1 = (((4'sd4)?(3'd1):(5'd14))?(~^(4'd14)):((2'd1)?(3'd1):(2'd1)));
  localparam [5:0] p2 = ((3'd4)?(3'd3):(3'd7));
  localparam signed [3:0] p3 = (3'sd0);
  localparam signed [4:0] p4 = ((4'sd1)>=(5'd8));
  localparam signed [5:0] p5 = (&(~^(-5'sd6)));
  localparam [3:0] p6 = (~^(2'd1));
  localparam [4:0] p7 = (!(~&{1{(^{2{{3{(&(-2'sd0))}}}})}}));
  localparam [5:0] p8 = (&(5'd0));
  localparam signed [3:0] p9 = (((4'd4)<<<(5'd23))<((3'sd2)==(5'd14)));
  localparam signed [4:0] p10 = (2'd2);
  localparam signed [5:0] p11 = (-{(5'd27)});
  localparam [3:0] p12 = ((!(|(((3'd2)<<<(-2'sd0))-((-3'sd0)&(3'sd1)))))<<(~|((6'd2 * (4'd7))||{1{((-4'sd5)===(4'd1))}})));
  localparam [4:0] p13 = {(!{((~(4'd13))!==((2'sd1)>(4'sd3))),{1{({(5'd12)}-((2'd3)==(3'd0)))}}})};
  localparam [5:0] p14 = (!(~(!(5'd25))));
  localparam signed [3:0] p15 = ((((3'd5)!==(3'sd3))|{1{(2'd1)}})?(((3'sd3)===(-2'sd1))^{2{(-4'sd6)}}):({4{(-4'sd7)}}^~((-5'sd4)?(4'sd5):(-5'sd15))));
  localparam signed [4:0] p16 = {(-4'sd5)};
  localparam signed [5:0] p17 = {2{(-(~^(&{4{(-4'sd2)}})))}};

  assign y0 = (~^($unsigned($signed(a4))?$signed({3{p6}}):$signed((a5?a5:a2))));
  assign y1 = {4{(^$signed(a0))}};
  assign y2 = (a2?b0:p0);
  assign y3 = (p13?p15:a3);
  assign y4 = (-3'sd2);
  assign y5 = {(-5'sd5)};
  assign y6 = (2'd1);
  assign y7 = $signed({({({a0})}>{{$signed(p17)}}),$unsigned({($signed(p0)<=(p12^~p15)),$signed({b5,p16})})});
  assign y8 = ((((-4'sd3)<=(p11?p9:p13))|(5'd27))-(5'sd7));
  assign y9 = (+((!(a5<<a2))>(2'sd1)));
  assign y10 = {{{({a3,a1})},(!(~$unsigned((|a0)))),$signed($unsigned((|{b5,b0})))}};
  assign y11 = (~^(-5'sd3));
  assign y12 = (-5'sd13);
  assign y13 = (+{{p10,p1,p2}});
  assign y14 = ((p2?p15:p3)?(3'd6):(p4?p7:p3));
  assign y15 = ((-4'sd7)^{(p8?b5:a1),(~&a0),(p10)});
  assign y16 = ($unsigned(($signed((-2'sd1))!={2{(4'd0)}})));
  assign y17 = {1{(-2'sd0)}};
endmodule
