module expression_00770(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(~(!(4'sd2))));
  localparam [4:0] p1 = (~&(|(~(|((|(~&((!(3'sd2))<=((5'sd2)&&(3'sd3)))))|{(((5'd8)>>>(2'sd0))-{(2'd1),(2'd1),(3'd5)})})))));
  localparam [5:0] p2 = ((6'd2 * ((2'd0)>>(5'd12)))>=((3'd4)<<<((3'd1)&&(-2'sd0))));
  localparam signed [3:0] p3 = {(2'd2),(5'd13),(2'd1)};
  localparam signed [4:0] p4 = (&(4'd2 * ((2'd1)?(4'd11):(3'd7))));
  localparam signed [5:0] p5 = (~^{{({(&(2'sd0)),((-2'sd0)||(5'sd9))}>>>(!(((4'd7)<<(-2'sd0))<((5'd30)!=(4'd6)))))}});
  localparam [3:0] p6 = ((4'd12)<<(3'd4));
  localparam [4:0] p7 = (((2'd0)>=(-5'sd10))|(~|(-4'sd6)));
  localparam [5:0] p8 = {2{{1{((-3'sd1)?(5'd3):(-3'sd1))}}}};
  localparam signed [3:0] p9 = ({1{{1{{1{((4'd12)&(-4'sd5))}}}}}}&({1{(-4'sd1)}}+((2'd2)&(2'd2))));
  localparam signed [4:0] p10 = (3'd7);
  localparam signed [5:0] p11 = {4{(2'sd1)}};
  localparam [3:0] p12 = {{4{{(4'd2)}}},(!(~&{(5'sd0),(5'sd8),(3'sd1)}))};
  localparam [4:0] p13 = (-(5'd25));
  localparam [5:0] p14 = ((((5'd31)>=(4'd15))>((-4'sd7)^(5'sd15)))>=(((5'sd13)<<(2'd2))!=((3'd3)||(2'd2))));
  localparam signed [3:0] p15 = ((^(~^{1{(4'd15)}}))+{2{((-5'sd2)||(-3'sd3))}});
  localparam signed [4:0] p16 = {3{{(3'd4),(5'd5),(-5'sd8)}}};
  localparam signed [5:0] p17 = (3'sd0);

  assign y0 = $unsigned(((-((p1?a2:p4)>=(4'sd0)))!=$unsigned((&((&(p15&p10))<<<(a2===b3))))));
  assign y1 = ((+((-3'sd0)<<<{(~|b5)}))!==(~(5'd13)));
  assign y2 = (~|$unsigned((~(~&({3{(p5)}}>(~^(3'd5)))))));
  assign y3 = {2{(a1?b0:p17)}};
  assign y4 = $unsigned($signed(p1));
  assign y5 = (({{a2,a3}}&{(b3===b0),(a5)})<=(({{(p3),{a1},{a0,b5}}})));
  assign y6 = ($unsigned(b5)<=(b5==p15));
  assign y7 = ((+(4'sd0))==(-5'sd10));
  assign y8 = (-2'sd0);
  assign y9 = {1{{3{(!a4)}}}};
  assign y10 = {2{((a2||a3)!=={3{a3}})}};
  assign y11 = ((-2'sd0)<=(a2?a2:a4));
  assign y12 = $unsigned(({$unsigned({(b4),{p9},(-3'sd0)})}<<{{p14,p15},((4'd13)),(p17<p8)}));
  assign y13 = ({3{(|b2)}});
  assign y14 = (^$unsigned((~$unsigned((-(-5'sd13))))));
  assign y15 = (~^(^(~|$unsigned((p11)))));
  assign y16 = ((((a1||p3)>=(p17!=b4))<((p11||p10)<<<(a0&&a2)))>=((b4^~p11)/p13));
  assign y17 = {b4,b2,a0};
endmodule
