module expression_00639(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd1)*(2'd1));
  localparam [4:0] p1 = (^(+(!{(-4'sd6),(-2'sd1)})));
  localparam [5:0] p2 = {{({(2'd0)}>=((3'd0)<(2'd2))),(((5'sd2)<<<(5'd30))!=((-4'sd0)>=(-3'sd1)))}};
  localparam signed [3:0] p3 = (-5'sd9);
  localparam signed [4:0] p4 = ((((5'd30)?(-5'sd3):(4'd0))?{(4'd3),(4'd8),(5'sd12)}:{(5'd9),(5'd16)})!==(((2'sd0)>>(5'd10))<<{((3'd3)?(5'd31):(3'd6))}));
  localparam signed [5:0] p5 = (~&(-2'sd1));
  localparam [3:0] p6 = (+(!{2{{3{(3'd4)}}}}));
  localparam [4:0] p7 = {4{({(2'd1),(3'd2),(3'sd2)}^~{(3'sd1),(3'sd1)})}};
  localparam [5:0] p8 = (-3'sd0);
  localparam signed [3:0] p9 = (^{2{(&(+(3'sd0)))}});
  localparam signed [4:0] p10 = (+(((~^(2'd3))+((-2'sd0)&&(3'sd2)))===(+{(5'sd3),(3'd4)})));
  localparam signed [5:0] p11 = {3{{4{(-4'sd5)}}}};
  localparam [3:0] p12 = (((4'd5)?(4'd3):(4'd14))>>(~(4'sd2)));
  localparam [4:0] p13 = (((-4'sd2)|(4'sd6))?((5'sd10)^(5'd19)):((3'sd2)+(-3'sd0)));
  localparam [5:0] p14 = ((&((2'd0)<(2'sd1)))&(~|((-5'sd15)^(3'd6))));
  localparam signed [3:0] p15 = {2{(~&{2{(6'd2 * (4'd13))}})}};
  localparam signed [4:0] p16 = ((5'd25)?(2'd2):(-3'sd3));
  localparam signed [5:0] p17 = ((((4'd15)^~(4'd12))?((4'd1)^~(-5'sd14)):((5'sd4)?(-3'sd1):(2'd0)))?(((5'd6)^~(5'd22))!==((5'd25)?(4'd15):(4'd4))):(((-3'sd2)||(2'sd1))?((-2'sd1)?(3'sd0):(4'd7)):((3'd0)^(5'd10))));

  assign y0 = ((p13>=p0)?$unsigned((b0?a4:p2)):(-(&a0)));
  assign y1 = ((5'd29)&&(2'd3));
  assign y2 = ((4'd2 * (p14==p14))||$unsigned(($unsigned((p3?p0:p3))||$unsigned({a4,p14}))));
  assign y3 = {(&p1),(^p17),(~|p11)};
  assign y4 = (4'sd0);
  assign y5 = (({a3,a1,b0}+(b1+a2))!==((a0-a5)|(a2^~a1)));
  assign y6 = ((3'd0)?(a4!=a4):(~(~|b4)));
  assign y7 = $unsigned(((-3'sd0)!==((b3|a1)<<(b4||b1))));
  assign y8 = ((-3'sd2)&((^(b3!=a2))!==$signed((!(^a3)))));
  assign y9 = {4{p9}};
  assign y10 = $signed(p16);
  assign y11 = {1{({{1{((+a5)?(p2?b5:b5):$unsigned(a4))}}}<<<(&{4{(p12<=b5)}}))}};
  assign y12 = {3{a5}};
  assign y13 = {1{{1{((|{3{a2}})?$signed((+{4{b3}})):({1{b4}}>(!p16)))}}}};
  assign y14 = (a1&&b1);
  assign y15 = (($unsigned((a3-a3))!==(b2&b1))>>(5'd7));
  assign y16 = (b0?b2:a1);
  assign y17 = $unsigned((6'd2 * a2));
endmodule
