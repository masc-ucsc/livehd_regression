module expression_00675(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(-2'sd1),(3'd3),(-3'sd1)}?((3'sd2)?(5'd3):(4'sd3)):{(4'd11),(2'd1)});
  localparam [4:0] p1 = ((-4'sd1)||({2{(5'd19)}}|{4{(-2'sd0)}}));
  localparam [5:0] p2 = ({2{((3'd6)&(-4'sd1))}}<({(-5'sd9)}?{2{(3'sd3)}}:(3'd4)));
  localparam signed [3:0] p3 = ({2{(((-5'sd8)|(2'd3))!==(|(-3'sd1)))}}^({4{(-2'sd0)}}<(((2'd3)&(4'sd1))<={1{(4'd3)}})));
  localparam signed [4:0] p4 = {3{(-5'sd0)}};
  localparam signed [5:0] p5 = (3'd5);
  localparam [3:0] p6 = (~|((4'sd4)<<<(2'd0)));
  localparam [4:0] p7 = ((5'd2 * (5'd2 * (5'd20)))>>>(((3'sd3)>(3'd1))&((4'sd6)<(4'sd5))));
  localparam [5:0] p8 = ((5'sd14)&(5'd19));
  localparam signed [3:0] p9 = (!(-5'sd3));
  localparam signed [4:0] p10 = (((5'd3)||(4'sd6))>>{1{(4'sd7)}});
  localparam signed [5:0] p11 = (~|((-3'sd0)&(-4'sd3)));
  localparam [3:0] p12 = (~^(|(2'd0)));
  localparam [4:0] p13 = (-((|(((4'd12)<<<(-4'sd7))^((2'd2)>(2'd3))))||(|(!((2'd3)&((3'd1)^~(-4'sd6)))))));
  localparam [5:0] p14 = {4{((-5'sd13)>>>(5'd15))}};
  localparam signed [3:0] p15 = (~&(3'd6));
  localparam signed [4:0] p16 = (~(2'd2));
  localparam signed [5:0] p17 = ((!(((4'sd0)<<<(-2'sd0))<=(|(-3'sd2))))&&{(5'd14),(&{(+(-2'sd0))})});

  assign y0 = {2{p11}};
  assign y1 = (+(b1|p2));
  assign y2 = (($signed((~(b5<<b5))))>>({4{b4}}+(a1^~p5)));
  assign y3 = (((a0>a0)<=$signed(a2))^(^(a3?a2:b5)));
  assign y4 = ({((a4+a4)==={b4,a3,a4}),(3'd5)}>>>({2{(p15||b0)}}>>>({{3{b4}}})));
  assign y5 = {(+((a0?b4:a1))),(~|(&{a3,p7,p4})),((|b2)?$unsigned(a1):{a3,a4})};
  assign y6 = (~^(a1?b0:a0));
  assign y7 = (a0?p4:b4);
  assign y8 = (!(((b4^b1)!==(b3-a1))-(~^{2{(p9^~p4)}})));
  assign y9 = (~|(~^{{3{{1{p1}}}},((p17?p7:p13)^(b5!==b0))}));
  assign y10 = {((|(a4?p17:p2))<<<$signed((+{1{p8}})))};
  assign y11 = ({3{(b1?a2:b3)}}!={3{(b4^~a3)}});
  assign y12 = ((-2'sd0)/p6);
  assign y13 = (~^(-2'sd1));
  assign y14 = ((b5?p14:b3)?((4'd2 * p2)>=(p12<<p16)):((p12%p0)>=(p13?b3:p13)));
  assign y15 = ({3{b0}}>=(p16));
  assign y16 = (~^(({4{a3}}?(|{a3,p13,b2}):{p10,p5,a2})|((b3?a0:b3)>=(~^{1{(b1<<b3)}}))));
  assign y17 = ({(a3?a0:a5),({2{a1}}<<<(b2||b4))}!=={1{({2{b3}}^{b4,b5})}});
endmodule
