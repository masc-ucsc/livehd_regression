module expression_00745(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-4'sd1)?(5'sd2):(2'sd1))^~((4'd15)?(4'sd6):(5'd22)));
  localparam [4:0] p1 = (((-2'sd0)*(5'sd7))<(+((-4'sd6)&(4'd13))));
  localparam [5:0] p2 = (((2'd2)?(-3'sd3):(-4'sd2))?{(-4'sd2),(-5'sd8),(5'sd13)}:{1{(5'd0)}});
  localparam signed [3:0] p3 = ({3{(4'd11)}}?((-5'sd11)<<<(-2'sd1)):{4{(4'sd5)}});
  localparam signed [4:0] p4 = ((2'd2)||(2'sd1));
  localparam signed [5:0] p5 = (5'd15);
  localparam [3:0] p6 = ({2{((4'sd7)?(-3'sd2):(4'd13))}}===(((2'sd1)==(4'd8))===((-5'sd3)+(-4'sd1))));
  localparam [4:0] p7 = ((4'd14)?(2'd2):(-2'sd1));
  localparam [5:0] p8 = {((3'd5)?(2'd0):(4'd11)),((4'd0)?(3'd7):(-4'sd2)),((3'd1)<<<(3'd1))};
  localparam signed [3:0] p9 = {3{{(~^{1{(2'd1)}})}}};
  localparam signed [4:0] p10 = {2{{(5'd23),(4'sd2),(5'd13)}}};
  localparam signed [5:0] p11 = (((-2'sd0)>(5'd5))%(5'd14));
  localparam [3:0] p12 = (~^(^(~&(2'sd0))));
  localparam [4:0] p13 = ({((5'd6)^~(2'sd1)),{(4'd3),(4'd10)}}<=({(2'd0),(-3'sd0)}?((3'd3)<<<(2'd0)):(4'd2 * (4'd9))));
  localparam [5:0] p14 = {1{({3{{3{(3'd6)}}}}>>(((3'd5)|(2'd3))^((5'd30)&&(2'sd1))))}};
  localparam signed [3:0] p15 = ({1{{1{((~&{3{(5'sd3)}})-{4{(4'sd7)}})}}}}==((5'd2 * (^(3'd3)))>=({2{(5'sd13)}}==(^(4'sd2)))));
  localparam signed [4:0] p16 = (5'sd13);
  localparam signed [5:0] p17 = (4'd0);

  assign y0 = {4{((b5||a5)!==(a0&&b2))}};
  assign y1 = {2{((~^$signed((b4==p11)))!={4{p10}})}};
  assign y2 = (a3!==a4);
  assign y3 = $signed({(p17?p17:p15),(p16?p9:b1),(p8<p11)});
  assign y4 = ((b5-p8)^~(5'd23));
  assign y5 = $signed((-3'sd0));
  assign y6 = (~^(&((5'sd13))));
  assign y7 = (((b4>>>b2)?(~^(~^p9)):(4'sd6))+{(p15?p4:p7),{b3,p1},(5'sd7)});
  assign y8 = ((^((a2?b1:p12)+(p7<<<b2)))?((p5?p0:p17)?(-5'sd1):(p6<=p14)):({p2,b0}||{p10,p14,a5}));
  assign y9 = (!(({p1,p7}<<<(p0<p6))<((a5|b2)!==(a5&&a5))));
  assign y10 = (6'd2 * (p8>p0));
  assign y11 = (4'd4);
  assign y12 = (^(~^(~^(~(((a2!=b0)>>(p16&&a4))-(~|(b1>>b2)))))));
  assign y13 = ((~(~a2))%p11);
  assign y14 = {3{((a4&a5)!=(p13||b5))}};
  assign y15 = ((-5'sd8)||{(2'sd0),{p4,a0},(-5'sd14)});
  assign y16 = {(~|(~&(^a5))),(!(!{b4,p0,a2})),(|{a1,a0})};
  assign y17 = (5'd20);
endmodule
