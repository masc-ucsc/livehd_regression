module expression_00444(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{2{(-3'sd2)}}}};
  localparam [4:0] p1 = (-(4'sd6));
  localparam [5:0] p2 = {3{((5'sd4)===(3'd1))}};
  localparam signed [3:0] p3 = (+(4'd1));
  localparam signed [4:0] p4 = {1{((((5'd2)&(3'sd3))!=={1{(3'd0)}})&(((5'd23)<=(5'd9))&{(4'd6),(5'sd0),(5'd8)}))}};
  localparam signed [5:0] p5 = ((!(-{((2'd3)!=(2'sd0))}))>>>{(|(-4'sd6)),((4'd1)==(3'd6)),((2'sd1)==(2'd3))});
  localparam [3:0] p6 = (((4'sd4)>=(3'd4))-((4'sd7)||(4'd3)));
  localparam [4:0] p7 = ((-3'sd2)>>(-3'sd3));
  localparam [5:0] p8 = {((3'd0)<=(5'd27)),((-5'sd6)|(3'sd2)),((-2'sd1)<(5'd1))};
  localparam signed [3:0] p9 = (((3'sd2)!==(5'd21))?((4'sd3)?(3'd5):(5'sd14)):(4'd2));
  localparam signed [4:0] p10 = (-{(((-3'sd3)+(2'sd0))>>((3'd6)<<<(2'd0))),(~^(|{(-4'sd1)})),{2{(|(4'd5))}}});
  localparam signed [5:0] p11 = ((((4'd0)?(5'sd11):(5'sd5))<=((-3'sd2)==(-5'sd9)))==(((5'sd8)>>(4'sd6))?((5'sd8)?(4'd3):(-3'sd2)):((-5'sd7)==(4'sd7))));
  localparam [3:0] p12 = ((2'sd0)-(((5'sd6)==(5'd22))^~((3'd6)+(2'd1))));
  localparam [4:0] p13 = ((+((-(2'd3))>=((3'd7)%(5'sd14))))>>>((~((2'sd1)>(5'sd14)))||(~&(!(3'sd3)))));
  localparam [5:0] p14 = ((5'sd7)-(3'sd1));
  localparam signed [3:0] p15 = {(-{1{(~^{2{(^(~((-5'sd14)?(5'd0):(-4'sd2))))}})}})};
  localparam signed [4:0] p16 = (2'd2);
  localparam signed [5:0] p17 = {{2{((5'd14)&&(5'd7))}}};

  assign y0 = {(2'd2),(2'd1),{4{a3}}};
  assign y1 = (({{a4}}==(b0!=a4))^~{(a4===b4),(a0!==b5)});
  assign y2 = (((~^(5'd5))<(+((p2>>p13)^~{p2,p15,p0})))&((~^(~(|(p2>>>p17))))&&{(+(p2<<p16))}));
  assign y3 = {{(&(!(~p10))),(~{p2,p4})},(&{(~{b2}),(|{p4})})};
  assign y4 = ((-2'sd0)-((2'd1)<(p14>b1)));
  assign y5 = (~{4{(b5?b0:a2)}});
  assign y6 = ((a2-b2)-(a2&p2));
  assign y7 = (|{1{($unsigned((($unsigned(a5)<=(p0>>>p1))))<<{4{{b0,a3,a4}}})}});
  assign y8 = ((^(p17?a4:p10))<<(^(p16?p2:p9)));
  assign y9 = (6'd2 * a2);
  assign y10 = (!(&a1));
  assign y11 = {4{b2}};
  assign y12 = ((3'd0)&(+{p3}));
  assign y13 = ({(-5'sd12)}>=({(b3&p15)}&$unsigned((b5|p15))));
  assign y14 = {1{(|((p9+b5)>=(~|(^b5))))}};
  assign y15 = (((p2||a0)&(p16%p4))-(3'sd0));
  assign y16 = {(4'd0),{(3'd6)},(4'd5)};
  assign y17 = {{{p16,p8},(6'd2 * p12),{4{p5}}}};
endmodule
