module expression_00619(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({(4'd12),(4'd5)}<=(~^(-2'sd1)))<=((~^(-5'sd13))>>{(4'sd0),(3'sd3)}));
  localparam [4:0] p1 = (~^{(((3'sd0)!==(4'd15))&&{(3'd0),(4'd13)}),({(-5'sd13),(-3'sd0)}&(~|(5'd4))),{((-2'sd0)===(4'd7)),{(5'd14)}}});
  localparam [5:0] p2 = ((((3'd2)^~(5'd30))<<{4{(-2'sd1)}})!=={3{(3'sd0)}});
  localparam signed [3:0] p3 = {((!(-5'sd8))<{(5'd16)}),{((2'd1)-(-2'sd0)),(-3'sd1)}};
  localparam signed [4:0] p4 = {(|{4{(2'd3)}}),(((5'sd6)>>>(-4'sd1))!=(~|(-4'sd4))),(((2'd1)^~(-5'sd12))?((-2'sd0)|(3'd2)):((-4'sd6)?(3'd4):(4'd13)))};
  localparam signed [5:0] p5 = {(((3'd5)!==(5'sd15))>=((2'sd1)?(2'd3):(4'd12))),(5'sd12),((3'd6)?{(3'sd3),(-5'sd4),(4'sd5)}:((4'sd4)>>(2'sd0)))};
  localparam [3:0] p6 = (&(!{(2'd0),(-3'sd0),(5'd19)}));
  localparam [4:0] p7 = (((2'd3)?(2'd3):(2'd2))?(3'sd2):(~{2{(3'd2)}}));
  localparam [5:0] p8 = ((5'd3)&(-2'sd0));
  localparam signed [3:0] p9 = ((((-5'sd7)>>>(2'd0))<=((-2'sd1)>(3'd7)))!=={1{(4'd14)}});
  localparam signed [4:0] p10 = (5'd3);
  localparam signed [5:0] p11 = (3'd7);
  localparam [3:0] p12 = {(5'sd15),(5'sd14)};
  localparam [4:0] p13 = {1{{3{(!(+{3{(2'sd0)}}))}}}};
  localparam [5:0] p14 = {(((3'd5)?(5'sd11):(-2'sd1))?((2'sd1)?(-3'sd3):(2'd0)):{(5'sd10)}),{1{{{2{(4'd7)}},((5'd29)?(2'sd0):(4'd5))}}}};
  localparam signed [3:0] p15 = (-5'sd13);
  localparam signed [4:0] p16 = ((+{(~|(4'd13))})!==({(-4'sd7),(5'd17)}^~{(3'd7),(3'd4),(-3'sd3)}));
  localparam signed [5:0] p17 = ((~((5'd9)?(2'd1):(3'd0)))>=((4'd1)+(5'd0)));

  assign y0 = (a0^p9);
  assign y1 = (^p10);
  assign y2 = (({1{(~(b3|a3))}}!==$signed((a5==b3)))!=(~|(4'sd4)));
  assign y3 = ($unsigned((p10?a0:p9))=={4{p7}});
  assign y4 = ((b5|p16));
  assign y5 = ((~^((&a4)?(|b4):(b1<<a4)))?(^({a3,a5}?(b4>>a5):(-p6))):(+{{b1,a4,a1},(a5>>>p4)}));
  assign y6 = ((-2'sd1)?(-4'sd3):((+p12)?{p2,p0}:(-3'sd2)));
  assign y7 = (2'd3);
  assign y8 = {$unsigned({{1{{b3,p9,a0}}},(6'd2 * b0),(b2<<<p4)}),({4{a4}}>>{{1{a3}},$unsigned(a5)})};
  assign y9 = ({(&a1),(b1-b5)}===(!{4{b4}}));
  assign y10 = (((p0>=p10)?(p15?p3:p12):(p16-p11))=={3{(p11+p3)}});
  assign y11 = (&(!(-$unsigned(({$signed((&(~a5)))})))));
  assign y12 = {({(p10?p8:p6),(p3<p4)}?((p14+p12)<(p9?p8:p17)):((a5?p17:p4)?(p9&&p2):(p12+p8)))};
  assign y13 = {((p0==p0)<(a4&&b3)),((p12>=b5)>>(+a1))};
  assign y14 = ((~&(4'd2 * p8))/p14);
  assign y15 = (((b4?b4:a4)>(b4?b0:p11))>>((b2*a0)?(b4<<<a4):(b4<<<p9)));
  assign y16 = (!{(~|(p9?b4:b4)),(p10?a2:p4),(6'd2 * (a0?b0:a1))});
  assign y17 = (^$signed({3{$unsigned({3{b0}})}}));
endmodule
