module expression_00073(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(-(((4'd4)-(-3'sd3))?(~|(-(-3'sd1))):(6'd2 * (4'd13)))));
  localparam [4:0] p1 = {3{((-5'sd15)+(5'd29))}};
  localparam [5:0] p2 = (5'd22);
  localparam signed [3:0] p3 = {((5'sd10)|(2'sd0)),{(2'sd1)}};
  localparam signed [4:0] p4 = (~^(~|(!(~(~^(-(~^(!(4'd12)))))))));
  localparam signed [5:0] p5 = {((2'sd1)|((5'sd5)===(4'sd1))),(((2'd2)?(-3'sd3):(-5'sd15))+(|(2'd2)))};
  localparam [3:0] p6 = (+(5'd22));
  localparam [4:0] p7 = (!({(2'sd1)}|((5'd9)!=(4'd4))));
  localparam [5:0] p8 = {(4'd14),{1{{(-3'sd1),(3'sd1),(5'd18)}}}};
  localparam signed [3:0] p9 = (2'd2);
  localparam signed [4:0] p10 = (-5'sd7);
  localparam signed [5:0] p11 = (((&(4'd11))&(4'd2 * (2'd2)))!==(((5'sd5)<<<(-4'sd3))===((5'd25)==(5'sd4))));
  localparam [3:0] p12 = (+(~^(!(~^(~&(~|(~&(-(~|(~|(~&{4{(4'd3)}})))))))))));
  localparam [4:0] p13 = (~^{4{(~^(+{1{(-3'sd2)}}))}});
  localparam [5:0] p14 = ((-5'sd14)^~(2'd1));
  localparam signed [3:0] p15 = (3'd4);
  localparam signed [4:0] p16 = ((((-3'sd3)?(3'd2):(3'sd3))|((-5'sd14)>(3'd5)))?({1{(5'sd10)}}==((2'd0)<<(5'd17))):(((-3'sd2)>>>(4'sd7))<=((5'd8)>(5'd12))));
  localparam signed [5:0] p17 = {{{2{{(5'd15)}}}},{{4{(5'sd11)}},{(-5'sd9),(4'd15),(3'd0)}}};

  assign y0 = ((~|(~&$unsigned((~$signed((2'd2)))))));
  assign y1 = ((~^{((5'sd10)),$signed((4'd0))})==({(2'd0),(-3'sd2),(b2)}!=(+(-3'sd2))));
  assign y2 = (((b3?p0:a2)-(-5'sd6))>>>((p6>>>a0)<<{2{a5}}));
  assign y3 = (+(^{{p2,p14},(-2'sd0)}));
  assign y4 = {({$unsigned((p0)),$unsigned({p14,p7,p16}),(p1<<<a4)}&&{{4{p10}},{{p8,p12,p11},(p17>=a2)}})};
  assign y5 = (p9?p6:a0);
  assign y6 = ((2'd0)<<{2{{2{(~^a1)}}}});
  assign y7 = $unsigned((^(2'sd1)));
  assign y8 = (p17-a0);
  assign y9 = (+(&{(~&{{4{p10}},{(&{1{{p1,p14,b3}}})},{{p9},{a1,p16},(~p16)}})}));
  assign y10 = (3'sd2);
  assign y11 = {4{(b0-p0)}};
  assign y12 = (4'd2 * (p6-p2));
  assign y13 = ({p4,p11}|(a4<=p12));
  assign y14 = {1{{2{(-3'sd0)}}}};
  assign y15 = ((2'd2)/p1);
  assign y16 = {{(6'd2 * b2),(4'd2 * p6),(p14|p17)},(({a5,a2,b3}<=(b0^~b0))!==((b4>>a1)&(b1^~b1)))};
  assign y17 = (~&(|{4{p13}}));
endmodule
