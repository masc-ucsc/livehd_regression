module expression_00373(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-5'sd13);
  localparam [4:0] p1 = (((-5'sd13)?(-5'sd13):(3'd0))?((3'd7)?(2'sd0):(2'sd1)):(((3'sd1)+(3'd5))<((2'd0)?(4'd15):(3'sd0))));
  localparam [5:0] p2 = ({{{(-3'sd2),(2'd2)}}}+((4'd2 * (5'd3))>>{2{(5'd14)}}));
  localparam signed [3:0] p3 = {((|(4'd8))<<(~&(5'd22))),(4'd1)};
  localparam signed [4:0] p4 = (|(~(((!(-2'sd0))?((3'd5)?(3'sd0):(2'd1)):(~(3'd6)))?(~^(!((-2'sd0)?(3'sd3):(-3'sd3)))):(((3'sd3)?(-2'sd0):(-2'sd0))?((-2'sd0)?(3'd2):(3'd1)):((2'sd0)?(-5'sd3):(5'd22))))));
  localparam signed [5:0] p5 = (4'd2 * ((3'd6)>>(4'd7)));
  localparam [3:0] p6 = ((&({1{(5'sd8)}}==((3'd5)?(-5'sd15):(3'd5))))?(((5'd14)>>>(-4'sd4))>(-2'sd1)):(4'd2 * (3'd4)));
  localparam [4:0] p7 = ({(6'd2 * (5'd19)),((4'd10)>(5'd16)),((2'sd1)<<(4'd4))}|{4{{(3'd6),(-4'sd4),(4'sd3)}}});
  localparam [5:0] p8 = (3'd4);
  localparam signed [3:0] p9 = (|{2{(~|(4'sd6))}});
  localparam signed [4:0] p10 = (^(-(4'd15)));
  localparam signed [5:0] p11 = {(2'd1)};
  localparam [3:0] p12 = ((((5'd24)>=(5'sd9))&(|(5'd4)))^((-(4'sd7))!==(4'd7)));
  localparam [4:0] p13 = ((2'd3)!=(3'd3));
  localparam [5:0] p14 = {2{{4{(3'd6)}}}};
  localparam signed [3:0] p15 = (((-5'sd6)?(-3'sd2):(-4'sd6))!=(+(2'sd1)));
  localparam signed [4:0] p16 = ((((3'sd0)?(4'd6):(2'd2))===((-3'sd1)<<(4'd14)))!=((!(5'd15))<(~&(4'd6))));
  localparam signed [5:0] p17 = (({(2'd2)}&((5'd28)<(-5'sd13)))^{((3'd0)>=(2'd0)),((-4'sd3)-(5'd0))});

  assign y0 = {2{{3{{2{a5}}}}}};
  assign y1 = {3{(p3<<b4)}};
  assign y2 = (($signed({(5'd2 * a2)})==(3'sd0))>>>({(p0==p11),(p11<<<p17)}==(5'd30)));
  assign y3 = {(a3>a5),{a2,a0,b4},(5'sd7)};
  assign y4 = (+{(|((|(^p15))>={p9,b5,a0}))});
  assign y5 = (a1?a5:a2);
  assign y6 = (3'd3);
  assign y7 = (4'd2 * (b1!==a2));
  assign y8 = ((((+(p15>>>p15)))^((p7&p5)<<<(p17+b4)))^~(((a2<<a1)!==(b4>>a4))<<(6'd2 * (|p6))));
  assign y9 = (5'sd3);
  assign y10 = ((~|((b3?b4:p11)<(p13&p2)))=={((p13?p7:p1)+{(p13<<<p3)})});
  assign y11 = (({(b0|a5),{4{b3}}})==={{{b5,a1,a0},(a0==b5)}});
  assign y12 = (~&((p4<a3)|{1{b0}}));
  assign y13 = $unsigned({2{$signed((!((5'd2 * p0)|(p9|a4))))}});
  assign y14 = (!((a3&b3)+(5'sd2)));
  assign y15 = ($unsigned(((b1===b4)?{2{p12}}:(2'd3))));
  assign y16 = ((^(+(p11?a0:p13)))?{3{(a1?a0:p13)}}:(|(3'd0)));
  assign y17 = ((-(-2'sd1))>((p15?p15:p6)?(b1&a3):(~&a0)));
endmodule
