module expression_00020(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(~|{3{(5'sd10)}})}};
  localparam [4:0] p1 = ({3{(4'd7)}}?{2{(5'd26)}}:((3'd4)?(4'd10):(4'd13)));
  localparam [5:0] p2 = ((((2'd0)?(2'd3):(3'd4))||((5'd20)?(5'd27):(3'd3)))?(((5'sd5)?(2'd0):(3'd4))+((5'sd5)?(5'sd9):(-3'sd1))):((-5'sd4)?(4'sd1):(5'd28)));
  localparam signed [3:0] p3 = (((2'd0)|(3'sd3))<<<(4'd2 * (5'd31)));
  localparam signed [4:0] p4 = (~(-3'sd3));
  localparam signed [5:0] p5 = ((+((-5'sd9)?(2'sd0):(5'd5)))?((^(3'sd3))?(^(5'd29)):((-4'sd0)?(5'sd9):(4'sd1))):(~|(^((-2'sd1)?(5'sd13):(5'sd15)))));
  localparam [3:0] p6 = (~&(~^{(^{(~^({(4'd11),(3'sd3),(4'sd1)}>(|(&(2'd2)))))})}));
  localparam [4:0] p7 = (((2'd1)?(5'sd12):(5'd23))?((-5'sd12)-(4'd13)):((2'd3)==(3'd7)));
  localparam [5:0] p8 = (-(~|(|(~(({4{(5'd10)}}<<{1{(4'd3)}})+(|{(-5'sd6),(-2'sd1),(-5'sd8)}))))));
  localparam signed [3:0] p9 = (~{({{(-3'sd0),(4'd11),(4'd11)}}<{(3'd0),(5'd4),(3'd2)}),(((2'sd1)^(5'd3))&&{(3'sd0),(5'sd13),(3'sd3)})});
  localparam signed [4:0] p10 = (~^(!(&{3{{1{(5'd18)}}}})));
  localparam signed [5:0] p11 = ((|{(&(2'd3))})>>>{(~&(4'sd1)),(!(-2'sd1))});
  localparam [3:0] p12 = (((3'd1)?(2'sd0):(-4'sd6))>>((4'd1)?(3'sd0):(2'd1)));
  localparam [4:0] p13 = ((-4'sd6)===(2'd2));
  localparam [5:0] p14 = (4'd10);
  localparam signed [3:0] p15 = {(!((-3'sd1)?(5'd2):(5'sd11))),((3'sd0)?(5'd10):(2'sd0)),((3'd0)?(4'd1):(-3'sd3))};
  localparam signed [4:0] p16 = (|((-2'sd0)>(-3'sd2)));
  localparam signed [5:0] p17 = {((-3'sd0)?(2'd2):(4'sd0))};

  assign y0 = {1{{(-4'sd3),({p15,a1,p16}-{1{p2}}),({p6}<={p16,a3})}}};
  assign y1 = (((p8&a5)+(+b4))?{4{p4}}:(p12?a0:p1));
  assign y2 = ((!(5'd15)));
  assign y3 = {4{{1{{p17,b4}}}}};
  assign y4 = {(3'd0),({a1}?{b3,a4}:(5'sd4))};
  assign y5 = (((!b3)?(p1?p10:b5):(p13?a0:a3))?((a2^b5)&&(b0<<a1)):(~&(|(p7*a3))));
  assign y6 = (~&((~&(b5>>p16))^(^(b0^~b3))));
  assign y7 = ($signed($signed((3'd3))));
  assign y8 = (~($signed($signed(((~|p16)?(p16?p8:p10):(p0?p7:p8))))^~((((p6?p15:p14)?$unsigned(p16):(-p7))))));
  assign y9 = (((b2<p2)?{1{a0}}:(p17^~p9))?{4{(p1!=p7)}}:((p13^a3)?(p6?b3:b2):(p6?p14:a4)));
  assign y10 = (|(~(((a0>b5)&(a4?b2:a1))!==(~^(a2==a4)))));
  assign y11 = (5'd4);
  assign y12 = ({b3,a3,a4}=={b0});
  assign y13 = (4'd13);
  assign y14 = (^(^(+(|(&((^(+(a5|a4)))!=((~b3)!==(~a0))))))));
  assign y15 = ((b5!==b3)?(a0<=p17):(b3/a0));
  assign y16 = ((({4{p11}}==((-2'sd0))))?{4{(3'sd3)}}:($unsigned((b0!==a0))^~(4'sd2)));
  assign y17 = (^b1);
endmodule
