module expression_00056(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{{4{(3'd0)}}});
  localparam [4:0] p1 = (((4'd9)-(2'd2))?(-2'sd1):(3'sd1));
  localparam [5:0] p2 = {{(-5'sd2),(3'sd2)},((-5'sd5)&(2'sd1))};
  localparam signed [3:0] p3 = ((-4'sd4)&(4'd15));
  localparam signed [4:0] p4 = ((!(-3'sd2))>=((4'd9)?(-4'sd5):(4'd12)));
  localparam signed [5:0] p5 = (((2'd3)<(3'sd3))-(2'sd1));
  localparam [3:0] p6 = ((((5'd11)-(5'd11))>((-2'sd0)?(-2'sd0):(2'sd1)))?((5'd21)?(5'sd4):(3'sd1)):((4'sd3)?(2'd0):(2'd3)));
  localparam [4:0] p7 = (((3'sd1)!=(4'd6))%(3'sd0));
  localparam [5:0] p8 = {(4'sd6),(-2'sd0),(4'sd1)};
  localparam signed [3:0] p9 = ((-5'sd1)?(5'sd5):(2'd2));
  localparam signed [4:0] p10 = (-3'sd0);
  localparam signed [5:0] p11 = ({(-3'sd0),(3'd4)}?((2'd0)?(2'd0):(5'd0)):((-2'sd1)?(2'd3):(2'sd0)));
  localparam [3:0] p12 = (2'sd0);
  localparam [4:0] p13 = ((3'sd2)&&(((3'd0)^(-5'sd0))?{1{(3'sd0)}}:(-5'sd2)));
  localparam [5:0] p14 = (~(((^(2'd0))<<((2'd3)^(-5'sd3)))^((~(4'd13))&&((2'd1)!=(3'd7)))));
  localparam signed [3:0] p15 = (((&(6'd2 * (5'd31)))+(~^{(-4'sd4)}))!=(((-4'sd0)^~(-3'sd1))<<<(~^(3'd2))));
  localparam signed [4:0] p16 = (((2'sd1)?(4'sd5):(-3'sd2))?{(4'd4),(-3'sd0),(5'sd9)}:(|{(3'sd3)}));
  localparam signed [5:0] p17 = {(({((3'd6)|(-2'sd1))}>>((4'd0)||(-3'sd2)))!==(((5'd24)&&(2'sd0))>((2'd1)==(5'd26))))};

  assign y0 = (a2?p2:p2);
  assign y1 = (p3?p16:b3);
  assign y2 = (|{4{(!{{4{p5}},{2{a4}}})}});
  assign y3 = ({4{p8}}?((b1<b0)===(a2?b3:b4)):((b1?p3:p6)?(~&p11):{p3,p15,p6}));
  assign y4 = (({3{a5}}^((a0^b1)!={2{p7}}))^(({1{a0}}==(b0&a1))===({2{a5}}&(b4!==b1))));
  assign y5 = (~|(~(a1^~p6)));
  assign y6 = ({(~&(^a3)),{3{a1}}}!=(~(~&((4'd2 * b0)^~(p8||p7)))));
  assign y7 = (3'sd0);
  assign y8 = (^{4{(p13<=p10)}});
  assign y9 = ({2{{2{b2}}}}|{2{{b5,a4,b5}}});
  assign y10 = (a5?p15:p13);
  assign y11 = ((~|{2{b5}})==={2{a4}});
  assign y12 = {3{{2{(a4>>>b5)}}}};
  assign y13 = (~($unsigned((b1?p4:p7))?(p8?a4:a1):(p2?a5:a5)));
  assign y14 = (((-(~^p3))|(p11?p9:p14))<<$signed(((a0?p2:a0)!=(|p16))));
  assign y15 = ((a0*a1)*(~&(-4'sd5)));
  assign y16 = (((({4{b3}}?(a3^~a4):$unsigned(a5))))>>{3{$unsigned({3{b5}})}});
  assign y17 = $signed(((6'd2 * (~^(b1===a1)))));
endmodule
