module expression_00004(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(((2'sd1)?(-2'sd0):(5'sd10))?(^(+(-5'sd6))):(+(-(3'd7)))));
  localparam [4:0] p1 = (|({(4'd10),(-3'sd0),(-3'sd0)}?{(-(2'd3)),{(2'd3)}}:((-(3'sd1))||{(2'd2),(2'd1),(3'd6)})));
  localparam [5:0] p2 = (((5'sd1)?(3'd0):(5'd19))?((-5'sd14)?(4'd11):(4'd11)):((-4'sd7)^~(3'd0)));
  localparam signed [3:0] p3 = (2'sd0);
  localparam signed [4:0] p4 = (~(-5'sd15));
  localparam signed [5:0] p5 = (4'd2 * {(4'd3),(2'd2)});
  localparam [3:0] p6 = (((2'sd1)%(5'd1))>>((5'd7)?(4'd9):(4'd13)));
  localparam [4:0] p7 = {2{(((3'd3)||(-3'sd3))||{(4'd7),(4'd7)})}};
  localparam [5:0] p8 = {(((4'd7)?(5'd31):(2'd1))?{(&(5'sd1))}:{(4'sd1),(3'd6),(5'sd2)})};
  localparam signed [3:0] p9 = (!(4'd6));
  localparam signed [4:0] p10 = ({(4'sd0),(3'd5),(+(-3'sd0))}<<<(((4'sd0)<(3'd5))|(~|(4'd9))));
  localparam signed [5:0] p11 = {{(4'd14),(-5'sd8)}};
  localparam [3:0] p12 = (((!(5'd2))?(~|(-3'sd1)):(+(2'sd1)))?{(|(3'sd0)),((3'd2)<<<(4'd6)),((-3'sd3)>(-4'sd4))}:((|(-2'sd1))-((2'sd0)&(5'd10))));
  localparam [4:0] p13 = (-{3{(4'd0)}});
  localparam [5:0] p14 = ((((4'sd0)<(4'd9))&(-3'sd2))+(~(2'sd1)));
  localparam signed [3:0] p15 = (!{(&(3'd0)),(+(4'd12)),((-4'sd1)?(5'd17):(5'd17))});
  localparam signed [4:0] p16 = ((4'd2 * ((5'd9)>(3'd2)))?(-3'sd3):((4'd9)?(5'sd15):(-2'sd1)));
  localparam signed [5:0] p17 = {4{(&(5'sd9))}};

  assign y0 = (((~&$unsigned(p6))^~{p14,p15})<<<({a0,a3}!==(a5<<<a1)));
  assign y1 = ((5'd7)^~((4'sd1)?$unsigned(p17):(p9==b0)));
  assign y2 = {1{(((p17!=p16)?(p15?b2:b1):(b2?a2:b5))?{3{(~b2)}}:(~&(|{4{p0}})))}};
  assign y3 = (({4{a5}}!={2{(4'd2 * p12)}}));
  assign y4 = ((~&(^(p3&a3)))<=((|p15)<<(!a4)));
  assign y5 = (!{(-2'sd1),{(4'd8)}});
  assign y6 = (+(-3'sd0));
  assign y7 = {(|(b5)),(p7||p1),{1{(~|p14)}}};
  assign y8 = $unsigned(($unsigned(p12)));
  assign y9 = $signed((a2?a4:b1));
  assign y10 = (~&({(p13||a2)}>={p9,p14,p10}));
  assign y11 = {{{{$unsigned(p16),{p13,b2}},$signed({p13,a4}),{2{{2{p12}}}}}}};
  assign y12 = {3{(b3?p10:a1)}};
  assign y13 = {{3{(b3>>b1)}},{1{({4{a0}}?(p2?b2:p8):{4{p17}})}}};
  assign y14 = (-((a3&b3)||(3'sd2)));
  assign y15 = $signed((~((4'd8)>>$unsigned(((p11>>b5)>=(!b5))))));
  assign y16 = (2'd1);
  assign y17 = (3'sd3);
endmodule
