module expression_00521(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~((-4'sd1)?(3'd1):(3'd1)))?((5'sd15)===(5'd10)):((3'd6)^(3'd0)));
  localparam [4:0] p1 = {3{{3{(2'sd1)}}}};
  localparam [5:0] p2 = (&(~(4'd11)));
  localparam signed [3:0] p3 = ((5'sd9)>>>(-5'sd2));
  localparam signed [4:0] p4 = {4{{3{(2'd3)}}}};
  localparam signed [5:0] p5 = ({(+(+(6'd2 * (2'd2))))}=={{(~&((4'd11)||(5'd9)))}});
  localparam [3:0] p6 = (~&(~(|(3'sd0))));
  localparam [4:0] p7 = {1{((2'd1)+(-5'sd1))}};
  localparam [5:0] p8 = ((((5'd20)?(5'sd1):(2'd2))?((-3'sd0)?(3'd1):(-3'sd0)):((-4'sd5)?(3'sd0):(5'd14)))?(((-5'sd1)?(5'sd12):(5'sd14))?((2'd2)?(4'd5):(4'd5)):((5'sd3)?(5'd18):(4'sd6))):(((4'd2)?(-4'sd6):(4'sd3))?((4'd4)?(5'd29):(3'd2)):((5'sd6)?(-5'sd7):(-2'sd1))));
  localparam signed [3:0] p9 = (4'sd6);
  localparam signed [4:0] p10 = ((3'd0)^~(5'd15));
  localparam signed [5:0] p11 = (+(-5'sd4));
  localparam [3:0] p12 = (&(&(|(3'd2))));
  localparam [4:0] p13 = ((((-2'sd1)|(5'd22))<<((3'sd0)-(3'd7)))?(((-5'sd2)?(-3'sd1):(-4'sd1))||((-4'sd4)==(3'sd2))):(((2'd3)+(4'sd1))?((-4'sd6)<=(4'sd2)):((3'd2)>>(-5'sd11))));
  localparam [5:0] p14 = {4{(((3'd6)<(4'd8))&{1{(3'd7)}})}};
  localparam signed [3:0] p15 = (!{2{(((-5'sd11)<<(3'd1))=={2{(5'd14)}})}});
  localparam signed [4:0] p16 = (2'sd1);
  localparam signed [5:0] p17 = ((((5'sd15)*(5'sd11))<=((2'd3)|(-3'sd3)))!=(((5'd0)<(4'd9))||((2'd2)%(4'd9))));

  assign y0 = (((~&a5)^~(b2!==a3))!==(-$signed((~(b0^b1)))));
  assign y1 = ($unsigned(p3)/p0);
  assign y2 = (&{{(&{p16,p8,p9}),{2{{4{p0}}}}},({3{b1}}<<(-(a1!==b1)))});
  assign y3 = (~|(!(((&b4)<<<(~^a2))?(p12?b4:b2):((a4&b1)%a5))));
  assign y4 = {(~&(~&(2'sd1)))};
  assign y5 = {(a1^p4),(b1==a3)};
  assign y6 = {b5,b0};
  assign y7 = {$signed((2'd3))};
  assign y8 = (4'd4);
  assign y9 = ((($signed(({((a1?a5:b5)?{p14,a3}:(a4?p15:a0))})))<($unsigned((b0<b5))?$unsigned($unsigned(a2)):(p9?a0:a2))));
  assign y10 = (((b0?a1:a5)===(&(|a4)))==(^((a0?b3:a5)?(~|a4):(-b4))));
  assign y11 = (((5'd12)));
  assign y12 = (((p3?a4:b3)>>>(b5?p16:p7))-{4{$signed(b3)}});
  assign y13 = (p5&&p10);
  assign y14 = ({3{(p16?b2:b0)}}>>>{{3{a4}},((b2?a3:a0)-(p13>=b1))});
  assign y15 = (p13?p4:p4);
  assign y16 = ((p6?a0:b1)<(p12<=b5));
  assign y17 = (~{3{$unsigned((-3'sd3))}});
endmodule
