module expression_00940(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'sd5)>(5'd22))<<<(5'd2 * (5'd14)))!==(((3'd1)-(-3'sd0))&&((5'd19)==(2'd2))));
  localparam [4:0] p1 = (^(((-5'sd15)>>(3'd5))<(|(&(-2'sd0)))));
  localparam [5:0] p2 = {3{{{(-2'sd1),(5'd0),(4'sd5)},{(-4'sd3),(5'd9)}}}};
  localparam signed [3:0] p3 = (5'd2 * ((2'd2)<=(4'd1)));
  localparam signed [4:0] p4 = ((3'd7)-({(2'd2),(-4'sd6),(4'd3)}>>(-4'sd0)));
  localparam signed [5:0] p5 = {4{(3'd0)}};
  localparam [3:0] p6 = (-(((3'd4)?(3'd6):(2'd2))%(2'sd1)));
  localparam [4:0] p7 = ((&((5'sd5)<(3'd3)))<<(&(-(4'd8))));
  localparam [5:0] p8 = (((2'd3)?(2'sd1):(2'd2))?{(3'sd3),(2'd0),(2'd2)}:(2'd3));
  localparam signed [3:0] p9 = (~|(((4'sd4)>>((4'd13)===(-2'sd1)))?((4'd10)>(-(-2'sd1))):((6'd2 * (5'd17))?(5'd2 * (4'd14)):(^(3'd5)))));
  localparam signed [4:0] p10 = ((2'd0)^~(3'd0));
  localparam signed [5:0] p11 = (((3'd3)^~(3'sd0))||{(4'sd2),(4'sd2)});
  localparam [3:0] p12 = (((-2'sd1)!==(2'sd1))<=((3'd3)<<(-2'sd0)));
  localparam [4:0] p13 = ((|(4'd15))<<<{(-2'sd1),(4'd0),(3'd7)});
  localparam [5:0] p14 = (((4'd11)<(-4'sd4))<((5'sd7)||(-5'sd8)));
  localparam signed [3:0] p15 = ((4'd2 * (4'd0))/(5'sd8));
  localparam signed [4:0] p16 = (-(|((((-2'sd1)&(-2'sd0))||{(-3'sd3),(4'd14)})=={{(-4'sd0),(3'd4)},((-5'sd8)>=(2'sd1))})));
  localparam signed [5:0] p17 = {1{(&({2{(3'sd2)}}?(^((-4'sd0)?(4'sd6):(5'sd8))):((3'sd0)?(3'd2):(2'sd0))))}};

  assign y0 = {1{((p12?p7:p0)?{4{p3}}:(2'sd0))}};
  assign y1 = (^(!((^(p14?p2:p12))|(-{p3,a5,p12}))));
  assign y2 = (((p7<=p1)+(p15?a4:p11))?($unsigned({4{a3}})):(({1{(p2?p5:b5)}}||(p10?b3:p5))));
  assign y3 = (({a3}+{4{p15}})=={(~^b5),(a3!=a3)});
  assign y4 = (-(&(5'd18)));
  assign y5 = (3'd5);
  assign y6 = ((p2==a4)^(a2^p13));
  assign y7 = ((|b5)/p7);
  assign y8 = ({3{{p4,p12,p15}}}>{4{{b5,p12,p10}}});
  assign y9 = ((a2&&p0)+(b2>p6));
  assign y10 = (6'd2 * $unsigned((^a5)));
  assign y11 = (3'd5);
  assign y12 = (b5>>>p9);
  assign y13 = (~(~&b2));
  assign y14 = ((3'd5)^~(a1?b1:a0));
  assign y15 = (((a1?b0:b3)|(b2?a1:b3))<<<((b4==p13)?(a0^b4):(a5&&b3)));
  assign y16 = (((a5-a2)==(b3+a3))<(|{(p16==b2)}));
  assign y17 = (~&(^$signed((^{({{(-3'sd0)}}+({p2,a4}!=(-5'sd2))),((3'd0)==(4'd8))}))));
endmodule
