module expression_00211(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd7)?(4'd8):(4'd2))?((3'd2)?(-2'sd0):(-2'sd0)):((3'd5)?(4'sd1):(-3'sd2)));
  localparam [4:0] p1 = (^((~(3'd1))<=((2'd1)<=(-2'sd1))));
  localparam [5:0] p2 = (!(^(-4'sd0)));
  localparam signed [3:0] p3 = ({4{(5'd10)}}?{{1{((4'd10)?(-4'sd6):(3'd6))}}}:{1{(5'd2 * (4'd5))}});
  localparam signed [4:0] p4 = (((-2'sd0)?(2'd2):(5'd28))?((5'd20)-(2'sd0)):((-3'sd1)|(2'd0)));
  localparam signed [5:0] p5 = (((2'sd0)<<<(3'd5))/(5'sd8));
  localparam [3:0] p6 = ((-3'sd3)!=(2'd1));
  localparam [4:0] p7 = ({(4'sd1),(-4'sd5)}&((4'd14)+(2'sd1)));
  localparam [5:0] p8 = ((~^((5'd9)==(4'd6)))!=={3{(4'd1)}});
  localparam signed [3:0] p9 = (!(|{{3{(~|(2'sd0))}}}));
  localparam signed [4:0] p10 = (~((~^{({(5'd4),(5'd16),(4'sd4)}===(-3'sd0))})^~(-4'sd2)));
  localparam signed [5:0] p11 = (((+(2'd0))?(~&(-5'sd12)):(|(-3'sd1)))?(((5'd11)?(2'sd0):(4'sd4))?((3'd2)>=(-4'sd3)):((-3'sd1)?(2'sd0):(4'd9))):(+((3'sd0)?(2'sd0):(4'd12))));
  localparam [3:0] p12 = {2{(-3'sd1)}};
  localparam [4:0] p13 = ({2{((5'd19)?(3'd3):(2'd3))}}>>(((-4'sd1)?(3'sd1):(2'd1))?((5'sd10)&(3'd6)):{1{(3'sd1)}}));
  localparam [5:0] p14 = (~(((-4'sd1)<<(4'sd3))?(-3'sd1):((4'sd3)?(4'sd5):(-5'sd10))));
  localparam signed [3:0] p15 = (3'd3);
  localparam signed [4:0] p16 = (((4'd14)?(4'd0):(-5'sd0))?((-5'sd15)?(-5'sd0):(4'sd4)):{2{((3'sd2)?(4'd12):(5'd25))}});
  localparam signed [5:0] p17 = {(5'd30),(2'sd0),(-5'sd4)};

  assign y0 = ((p15?b1:b1)?(p16?p17:a2):(p16?p4:p15));
  assign y1 = (a1?b5:b3);
  assign y2 = {{(a2>>p1),(p16)}};
  assign y3 = (5'sd1);
  assign y4 = ((3'd7)!==(((b3&a1)>>>(a1>>a1))+((2'd2)&&{4{a4}})));
  assign y5 = (~^(5'd2 * (-(5'd30))));
  assign y6 = ((b3?p13:p7)?(-p11):(a2<b1));
  assign y7 = (~&(|(~|((&({2{p7}}||{4{b4}}))<<((^((~|p15)<<(p5?p4:b5))))))));
  assign y8 = ((3'sd0)^~(~^b4));
  assign y9 = (&$unsigned((p12<=p16)));
  assign y10 = (((b5==p5)|(a5!==a1))+({3{a2}}!==(b4!==b1)));
  assign y11 = (6'd2 * $unsigned((a3!==b4)));
  assign y12 = {3{{3{(-4'sd6)}}}};
  assign y13 = (((&(4'sd1))<=(b5?a4:b0))===((|(4'sd3))!==(a0?a5:b1)));
  assign y14 = (^{p9,a3});
  assign y15 = ((^a5)<<<(b5^~a0));
  assign y16 = (~{(~{{b2},(-b2)}),({a3,b2}==={a3,b0,a5})});
  assign y17 = {(p15?b3:b2),(p10?a1:a2),(a0?a4:a3)};
endmodule
