module expression_00047(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^(3'd1))?((-2'sd1)<=(-2'sd1)):((3'd1)!=(4'd9)));
  localparam [4:0] p1 = (^(|(~|(~|(+(~&(~&(&(-(~&(-5'sd7)))))))))));
  localparam [5:0] p2 = {{(5'd24),(-4'sd6),(4'sd5)},(~&{(5'sd0),(5'd17)}),(((3'd5)<=(4'sd2))!=((5'd25)|(3'd5)))};
  localparam signed [3:0] p3 = (~(~^(-3'sd3)));
  localparam signed [4:0] p4 = (({(+{(-2'sd0),(-5'sd12)})}&&((|(5'd25))<<<(!(4'd11))))>({(-5'sd7),(3'd4),(4'd1)}|(|(~^((-3'sd2)>(2'sd1))))));
  localparam signed [5:0] p5 = (!(!(&(&(2'sd1)))));
  localparam [3:0] p6 = {{{{1{{3{(-3'sd2)}}}}},{1{{{4{(5'sd14)}}}}}},{{({{1{(2'd2)}}}<=((3'd4)>>>(3'sd0)))}}};
  localparam [4:0] p7 = {3{{3{((2'd0)-(2'sd1))}}}};
  localparam [5:0] p8 = (|((((5'd12)>=(5'sd9))^(!((3'd1)||(5'sd4))))|((+(4'd2 * (4'd10)))||((2'd0)^~(-5'sd1)))));
  localparam signed [3:0] p9 = {4{(2'd2)}};
  localparam signed [4:0] p10 = ({(4'sd2),(5'sd8)}>>>(~&(4'd2 * (3'd6))));
  localparam signed [5:0] p11 = {(2'd3),(4'd12),(-5'sd5)};
  localparam [3:0] p12 = (5'd19);
  localparam [4:0] p13 = (!(3'd2));
  localparam [5:0] p14 = ((((3'd1)<=(2'sd1))===((4'sd2)?(-5'sd13):(4'sd3)))||(-5'sd5));
  localparam signed [3:0] p15 = ((2'sd1)?(4'd1):(4'sd2));
  localparam signed [4:0] p16 = {(4'd7),(3'd4),(4'd3)};
  localparam signed [5:0] p17 = ((-4'sd5)||((2'd2)?(-4'sd7):(5'd1)));

  assign y0 = (-3'sd3);
  assign y1 = (((b1?p17:b0)?(|p11):(p11>p11))?(~&(6'd2 * (p14==p0))):(~(5'd2 * (p12?p2:p6))));
  assign y2 = (&(+(~|(|(~^(^(~{1{({(^b4),(-a3),(b4?b2:b4)}!=({a0,b5,b3}-{3{b4}}))}})))))));
  assign y3 = ((~^b0));
  assign y4 = $unsigned((-($unsigned($unsigned(((!p7))))&((p2<=p1)==$unsigned(p1)))));
  assign y5 = (+{(~&b2),{a5,a3},{1{a1}}});
  assign y6 = ({1{{(5'd2 * a2)}}}?((~|p0)?{p0,p9}:{4{p16}}):{1{(+{2{b0}})}});
  assign y7 = ((((6'd2 * a2)!==(a0<a5))<<<((p6^~b0)==(a4/p14)))!=(((b3&&a1)^~(a4!=b4))!==((b1&a3)==(b0&b3))));
  assign y8 = ($unsigned(((p1?b0:p11)^{4{b2}}))<($signed((|((a2||a5)?(b3!=p3):(b2?b0:a0))))));
  assign y9 = (((4'sd4)&((4'sd1)*(a3!==a1)))<<(((3'sd1)<<(5'd21))-((b3^~a5)<(b1^~p14))));
  assign y10 = (2'd2);
  assign y11 = $unsigned({(!$signed((((p14||p0))>>>(a2^~p8))))});
  assign y12 = (~|(3'sd1));
  assign y13 = {2{((~&a0))}};
  assign y14 = {2{(p10?p6:p16)}};
  assign y15 = (((~|b2)&&(a3-b4))>={{2{b0}},(a3>p14)});
  assign y16 = ((b5-b2)/a1);
  assign y17 = ((((a1>>a0))!=={2{(a4<<b2)}})>>>(((^b1)>>(~^p8))-((~a2)<(6'd2 * p2))));
endmodule
