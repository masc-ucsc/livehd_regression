module expression_00510(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd13)<<<(5'd30))<<{4{(5'd16)}})>>>({4{(2'd2)}}<<{2{(-2'sd0)}}));
  localparam [4:0] p1 = (((3'd2)>((4'd12)^(4'd6)))?(((3'sd2)^~(3'd7))+((-3'sd0)==(3'sd2))):(((2'sd1)&&(4'd5))<<(5'sd4)));
  localparam [5:0] p2 = (-5'sd1);
  localparam signed [3:0] p3 = {{(4'd14),(5'd31)},{(5'd18),(2'sd0)}};
  localparam signed [4:0] p4 = (((4'sd5)?(4'sd5):(-3'sd0))?((5'd6)?(-3'sd2):(4'd7)):(3'd6));
  localparam signed [5:0] p5 = (~(3'sd2));
  localparam [3:0] p6 = {(6'd2 * {((5'd12)<<(4'd1))})};
  localparam [4:0] p7 = (5'd18);
  localparam [5:0] p8 = {((&(5'd8))?(-(5'd25)):(+(2'sd1))),(((4'sd5)?(4'd4):(5'd29))?((2'sd0)|(-5'sd5)):((3'd1)>=(5'sd12))),({(-4'sd5),(2'sd0)}&&{(2'sd1),(5'sd11),(-5'sd7)})};
  localparam signed [3:0] p9 = {(6'd2 * (3'd6)),((4'd8)?(3'd0):(3'sd1))};
  localparam signed [4:0] p10 = ((5'd9)?(3'sd0):(2'sd0));
  localparam signed [5:0] p11 = (2'd1);
  localparam [3:0] p12 = ((~{4{(5'd3)}})?(-((5'sd7)?(-3'sd0):(3'd3))):(|{4{(3'd5)}}));
  localparam [4:0] p13 = ((((2'sd0)?(-2'sd1):(5'd2))?(4'd6):{(4'd3),(5'd31),(5'd9)})?{(|(2'sd0)),{(-4'sd4),(-2'sd0),(3'd5)},{(5'd11),(3'd1),(3'd7)}}:(2'd0));
  localparam [5:0] p14 = (((-4'sd1)||(4'sd3))!==(+(~(-2'sd0))));
  localparam signed [3:0] p15 = {(&({({(5'sd10),(4'sd5),(4'sd1)}>={(5'd29),(-5'sd9),(2'd2)})}>>{{(-3'sd3)},{(-3'sd0),(-5'sd14),(-2'sd0)},(+(-5'sd10))}))};
  localparam signed [4:0] p16 = {4{(-(2'd1))}};
  localparam signed [5:0] p17 = ({3{((2'd3)+(4'd12))}}<=(((5'd20)!=(5'd22))?((5'sd9)<=(5'sd6)):(4'd2 * (4'd3))));

  assign y0 = (|(~({(a4?a3:a4),(2'd0)}<<{1{(~^{(2'd3),(a5===b5)})}})));
  assign y1 = ((p7?b0:p17)?{1{b1}}:(a3?a4:a3));
  assign y2 = (((p9<a0)?(a2===b3):(b2?a4:b3))!=$unsigned(((b4<=b1)?(~$signed(a2)):(-3'sd3))));
  assign y3 = ({4{(-2'sd0)}});
  assign y4 = (p14||a0);
  assign y5 = (((p2<<b2)|(p12^b3))<<(-((^(3'sd0))|(+(p16?b5:p17)))));
  assign y6 = ({{3{{2{a4}}}}});
  assign y7 = (|{({b1,a4}?{$signed(a3)}:(p6?a2:a1)),((p6?p17:p15)?(!(p12&&b3)):{b1,a4})});
  assign y8 = ((^((|(a2<<<a1))/p8))+(-((+(b3&b3))===((a5>a1)<(a5|a1)))));
  assign y9 = ({1{(3'sd0)}}?(4'sd0):((2'd1)?(3'd2):(p3>>>p2)));
  assign y10 = ((2'd0)&({1{a5}}>=(b5?b3:b1)));
  assign y11 = ($signed($signed(($signed((p4<p16))>=({3{p10}}==(p9>=a3))))));
  assign y12 = {1{{3{{3{b2}}}}}};
  assign y13 = (4'd9);
  assign y14 = ({b1,p4}?(a0?p2:b2):(b1?p11:p15));
  assign y15 = (($signed((4'd2 * a0))===($signed(a2)!==(a0^~b0)))>>($signed($unsigned((b4)))||$signed((a3<=a0))));
  assign y16 = (3'sd2);
  assign y17 = (~^(5'sd4));
endmodule
