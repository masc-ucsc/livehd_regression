module expression_00888(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd0)?(3'd3):(-2'sd0))?((3'd1)?(5'd24):(-2'sd0)):(+((4'sd6)^~(2'd3))));
  localparam [4:0] p1 = ((((4'd13)==((3'd4)!=(2'sd0)))<<<(^((-4'sd1)>>>(2'd1))))+{1{{1{((2'd1)||(-(~(2'd3))))}}}});
  localparam [5:0] p2 = ((5'd6)>>(-4'sd4));
  localparam signed [3:0] p3 = ((+((2'd1)?(3'd1):(5'd16)))?((-5'sd7)^(-2'sd1)):((-5'sd14)>>(2'sd1)));
  localparam signed [4:0] p4 = (((-3'sd2)<<(-3'sd2))==((5'sd1)*(3'd2)));
  localparam signed [5:0] p5 = {{(3'd0),(3'sd1),(5'd17)},(~^((2'sd1)<<<(3'sd1))),((5'd25)<<<(2'd2))};
  localparam [3:0] p6 = ({4{(-4'sd6)}}=={2{{1{(-4'sd1)}}}});
  localparam [4:0] p7 = (5'd18);
  localparam [5:0] p8 = ({((4'd4)?(-3'sd2):(5'sd5)),(5'd10),((3'sd3)?(5'd11):(4'd8))}?{{{(2'd1),(5'sd11)}}}:(~{(-4'sd2),(-4'sd0),(2'sd1)}));
  localparam signed [3:0] p9 = {4{(5'd2 * (5'd11))}};
  localparam signed [4:0] p10 = (~|(({(5'sd13)}>>>(~(-5'sd2)))+(&((+(4'sd0))^(+(4'd5))))));
  localparam signed [5:0] p11 = ((~&(4'd10))?((2'd2)<=(5'd25)):(5'd24));
  localparam [3:0] p12 = {2{{3{(3'sd0)}}}};
  localparam [4:0] p13 = (((5'd27)&(3'd4))!==(~^((-4'sd3)&&(-4'sd7))));
  localparam [5:0] p14 = (2'sd1);
  localparam signed [3:0] p15 = {3{{1{{1{((-3'sd3)^(-4'sd6))}}}}}};
  localparam signed [4:0] p16 = ((((-4'sd2)^(3'd5))<<<((5'd13)===(3'd5)))>((~(-2'sd1))||((4'sd4)<<<(2'd3))));
  localparam signed [5:0] p17 = (&{(5'sd9),(5'sd2)});

  assign y0 = {4{{3{p11}}}};
  assign y1 = (~&(~|(^(|($signed($signed((^(~|$signed(b0))))))))));
  assign y2 = (-4'sd5);
  assign y3 = ({(~^{(&(^(2'sd0))),(~({p17}?(-4'sd3):(-4'sd0)))})});
  assign y4 = (~^(a3/b2));
  assign y5 = $unsigned({{a1,b1,b3},{b1,p3}});
  assign y6 = (&(5'd28));
  assign y7 = (4'sd0);
  assign y8 = (((p0&p11)==(p8>>>p11))?((p10&&p11)):(p2?p6:a0));
  assign y9 = ({p0,a4,p1}<{(p12&b0),(a1?b1:p0)});
  assign y10 = {2{({1{(~(4'd4))}}>>({1{a5}}?(b3-b3):(~&p4)))}};
  assign y11 = {(|(({(~^{{$signed((~^p14))},$signed((~^(|a1)))})})))};
  assign y12 = {3{(5'd22)}};
  assign y13 = {2{{3{(b0&&a5)}}}};
  assign y14 = {1{(((((a1||p13))&$signed((p15<a2)))))}};
  assign y15 = (p17>a1);
  assign y16 = ((|((-a3)!==(a4>>>a5)))>>(~&(-((p9>a5)<<(b5===b2)))));
  assign y17 = {({{b0,p11},(^(+b4)),{b3,p16,a3}}&(({2{a2}}<<<(a2<<<a1))^((|b2)!==(~a4))))};
endmodule
