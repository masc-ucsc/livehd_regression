module expression_00094(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(|((4'd15)%(5'sd5))));
  localparam [4:0] p1 = ({(4'sd2),((-2'sd1)!==(-3'sd2))}!=(5'd10));
  localparam [5:0] p2 = (((3'd0)?(5'd30):(-2'sd0))<={2{((5'd21)?(4'd13):(4'd4))}});
  localparam signed [3:0] p3 = ((+(~(-(3'd6))))?(^((-5'sd11)?(-2'sd0):(4'd13))):(-((4'd7)?(3'd0):(3'd6))));
  localparam signed [4:0] p4 = (5'sd4);
  localparam signed [5:0] p5 = ((((2'd3)>>>(-4'sd3))&&((5'sd12)?(3'sd1):(5'd19)))||(3'd7));
  localparam [3:0] p6 = ((((2'd1)|(5'd3))&&((4'd13)+(-2'sd0)))<<((+(5'd4))>>(2'd3)));
  localparam [4:0] p7 = {3{(2'sd1)}};
  localparam [5:0] p8 = ({1{(4'd6)}}?((5'sd1)?(-5'sd9):(2'sd1)):((-5'sd0)?(-4'sd6):(-3'sd0)));
  localparam signed [3:0] p9 = ((((5'd12)>(-4'sd5))<=((3'd5)==(5'd30)))?(((4'd3)*(5'd27))>>>((-3'sd1)?(2'd2):(4'sd5))):(((4'd14)?(5'd11):(-5'sd9))<<((2'd1)<<<(3'd1))));
  localparam signed [4:0] p10 = (((-4'sd0)&&(4'd8))!=((3'sd2)^(4'd4)));
  localparam signed [5:0] p11 = ((~^{(~|(!(2'd1))),(^(|(3'd0)))})!==(^(~|(|(~{(5'sd15),(-3'sd1)})))));
  localparam [3:0] p12 = (((((-2'sd1)>(2'sd1))|((2'd1)+(5'd14)))>>(((-4'sd5)<(-3'sd0))===((5'd22)===(2'd1))))<=((((-3'sd0)+(4'sd1))+((5'd13)/(-5'sd1)))|(((5'd29)-(5'sd8))>>>((-3'sd1)*(3'd3)))));
  localparam [4:0] p13 = (!(~{(+{(4'd1),(-3'sd3),(4'd14)}),{(-4'sd0),(2'sd1)},(~|(|(5'sd1)))}));
  localparam [5:0] p14 = (~^(|(~^(-2'sd1))));
  localparam signed [3:0] p15 = {1{(5'sd8)}};
  localparam signed [4:0] p16 = ((4'd3)>=(((5'sd0)<=(5'sd13))<<<((2'sd0)||(3'd0))));
  localparam signed [5:0] p17 = {(((-3'sd1)^(4'sd0))?{(-4'sd6),(4'd3),(4'd10)}:(^(-5'sd10))),((|(4'd3))?{1{(2'sd1)}}:(^(5'sd1)))};

  assign y0 = {((a4!==a1)>>>{p16,b3,p7}),(-5'sd12)};
  assign y1 = (-5'sd14);
  assign y2 = {1{((b0===b1)?{1{(~|p13)}}:{2{a1}})}};
  assign y3 = (($unsigned((|b5))!==$unsigned({4{a5}}))+({4{p1}}>>(~(p13^a0))));
  assign y4 = {2{{{(p1?b4:p5),(b0?a5:b2)},(a2?p14:b5)}}};
  assign y5 = (((a1?b2:b0)-(b3?a5:b3))?{{(p8>p4)}}:$signed((a4?a5:a3)));
  assign y6 = ((-3'sd1)-(a2^p8));
  assign y7 = $unsigned({1{($unsigned((-{p17}))==(~|{{3{p10}}}))}});
  assign y8 = (((~|$signed(b3))/b5)>=((a2|b0)<<(-(b1))));
  assign y9 = ((5'd1)<<({p10,p8}||$unsigned((3'sd1))));
  assign y10 = (&(2'd2));
  assign y11 = $unsigned((({3{p5}}?{4{a4}}:{2{p5}})));
  assign y12 = {1{(^(+(~|{4{{1{({1{a4}})}}}})))}};
  assign y13 = {3{((^p9)?{3{p6}}:{1{p10}})}};
  assign y14 = {(-4'sd2),{(-3'sd1),$signed({b3,p4,p10})}};
  assign y15 = ((((3'sd1)!==(~&a4))<<(5'sd6))===(((4'd13)<<(2'sd1))>((~&b0)!==(b3-b1))));
  assign y16 = (((b0?p0:b2)>=(p14-b3))?((4'd2 * p6)+(p2?a5:p9)):((a5?p0:p1)/p4));
  assign y17 = {4{(a4?b1:a1)}};
endmodule
