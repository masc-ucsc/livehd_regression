module expression_00841(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd1)*(-2'sd0))>=((-3'sd2)>(4'd2)))<(((2'd3)*(2'd0))^((2'd0)<(3'd4))));
  localparam [4:0] p1 = ((4'd3)<(4'd11));
  localparam [5:0] p2 = (((2'sd1)===(2'd3))?((2'd0)<<<(3'd5)):((4'sd2)<=(4'sd3)));
  localparam signed [3:0] p3 = {1{({2{(-2'sd0)}}?((2'd2)?(-2'sd1):(3'sd0)):((5'd19)&&(4'd15)))}};
  localparam signed [4:0] p4 = {(2'd3)};
  localparam signed [5:0] p5 = (({4{(3'd4)}}||((3'sd1)!=(3'sd1)))>>{((3'd5)<<<(3'sd1)),((5'd30)^(-2'sd0))});
  localparam [3:0] p6 = (({(2'd0),(5'sd13)}-((3'd1)?(3'd3):(5'd20)))^~(((4'sd3)<<<(4'sd4))?((5'd12)+(2'sd0)):(~|(-4'sd2))));
  localparam [4:0] p7 = (-(&(~^(~^(~&(((~&(4'd8))>>(~&(5'sd0)))!=(|((-5'sd5)>(2'sd1)))))))));
  localparam [5:0] p8 = (^(-2'sd0));
  localparam signed [3:0] p9 = {2{{1{{4{{2{(4'd12)}}}}}}}};
  localparam signed [4:0] p10 = {2{(((5'sd0)>>>(-3'sd1))===((-5'sd13)<(3'd6)))}};
  localparam signed [5:0] p11 = (!{(-5'sd14),(3'sd2)});
  localparam [3:0] p12 = (^(4'd1));
  localparam [4:0] p13 = ((((4'd7)||(2'sd1))==={(3'sd0),(5'sd0)})?({(4'd0),(4'd11),(2'd3)}?{(5'd24),(-4'sd7),(3'sd2)}:((5'd0)&(4'd6))):{((4'sd2)>(3'sd2)),((4'sd0)?(-4'sd6):(2'd0))});
  localparam [5:0] p14 = ((-3'sd0)>>>(((3'sd3)<=(4'sd1))/(5'd22)));
  localparam signed [3:0] p15 = (|(5'd18));
  localparam signed [4:0] p16 = ((5'd23)<(-2'sd1));
  localparam signed [5:0] p17 = ((5'sd8)<=(2'd2));

  assign y0 = (~^{2{{1{(|p16)}}}});
  assign y1 = $unsigned((5'd20));
  assign y2 = {2{{3{b0}}}};
  assign y3 = (-4'sd4);
  assign y4 = {$signed(b4),{a0}};
  assign y5 = ($unsigned(p13)!=$signed(p14));
  assign y6 = (~(~|{2{(~|a2)}}));
  assign y7 = $signed($unsigned((((~&a4)+(b2&&a1)))));
  assign y8 = {{(a2?a1:b5),(a5?p6:b5),{b3}},((b0<=b0)+{(b1?b4:b0)}),((a5+b1)>(b5?p7:b2))};
  assign y9 = ($unsigned($unsigned($unsigned((p9))))?((a5)?(p11?a5:a0):(p16?a2:p17)):((p2?p17:a0)?(p10?p17:p3):(p6?b2:p17)));
  assign y10 = {p15};
  assign y11 = (~^p10);
  assign y12 = ((~|{4{a2}})?{4{a1}}:{4{b1}});
  assign y13 = (-5'sd10);
  assign y14 = ({(b5?b2:a5)}?(p6?p11:p10):{(a1?a1:a2)});
  assign y15 = ((b3?a5:a0)%b4);
  assign y16 = ((p4?p0:p4)^~(p15>b1));
  assign y17 = (({2{p11}}?(p2?p13:p5):(p0>>>p12))>=((4'd2 * p2)?{4{p13}}:{3{p16}}));
endmodule
