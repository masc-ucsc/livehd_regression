module expression_00860(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'sd2)>=(5'd22));
  localparam [4:0] p1 = (!(5'd22));
  localparam [5:0] p2 = ((4'd2 * (~|((4'd5)<(3'd5))))?(((-3'sd2)?(3'sd2):(5'd22))<<(~&(4'sd3))):(~((~|(-4'sd5))&&{(5'sd1)})));
  localparam signed [3:0] p3 = (4'd5);
  localparam signed [4:0] p4 = {1{((5'd8)<((-2'sd0)>>(2'd2)))}};
  localparam signed [5:0] p5 = (5'sd14);
  localparam [3:0] p6 = ((~((5'sd5)?(4'd5):(-2'sd1)))?{(~|(5'sd11))}:((3'sd0)?(-3'sd0):(4'd9)));
  localparam [4:0] p7 = ((4'd2 * ((3'd4)>>>(3'd2)))<{1{{3{(3'd3)}}}});
  localparam [5:0] p8 = (6'd2 * ((5'd15)||(3'd0)));
  localparam signed [3:0] p9 = {3{({4{(-2'sd0)}}>(5'd24))}};
  localparam signed [4:0] p10 = ((|({(5'sd14),(-5'sd0)}+((-3'sd3)===(-5'sd1))))>>({(2'd1)}?((3'sd0)<<<(3'sd0)):(+(2'd3))));
  localparam signed [5:0] p11 = (^(!(|(~|(5'd0)))));
  localparam [3:0] p12 = ((3'd5)||(-2'sd0));
  localparam [4:0] p13 = ({4{(5'd20)}}?(~(-3'sd3)):(6'd2 * (3'd7)));
  localparam [5:0] p14 = ((~|(|(~&(2'd1))))<(4'sd4));
  localparam signed [3:0] p15 = ((5'd8)?(-5'sd4):(5'sd11));
  localparam signed [4:0] p16 = (~|(+({4{(3'sd0)}}!=={2{(4'd9)}})));
  localparam signed [5:0] p17 = ({((2'd1)!==(3'd0)),(~&(5'd13)),{(5'sd7),(5'd7),(3'sd0)}}?(|(((3'd6)?(3'sd2):(4'd3))^~(+(4'sd0)))):((&(3'd1))!==(~(5'd29))));

  assign y0 = (({4{b2}})-((b5?b4:a0)^~(~^b2)));
  assign y1 = (5'sd8);
  assign y2 = (((~(|(!(p16<<b3))))!=(2'd0)));
  assign y3 = {1{(&p1)}};
  assign y4 = (~&$unsigned((-4'sd3)));
  assign y5 = (4'sd6);
  assign y6 = (2'sd0);
  assign y7 = (+((|($signed({a4,p11,b2})>=(p14^~a3)))));
  assign y8 = (|(!(-(4'd15))));
  assign y9 = {2{(p0!=p13)}};
  assign y10 = (-4'sd5);
  assign y11 = (((a5<<p14)^(&b4))?($unsigned(p7)<=$unsigned(a1)):(~((a2|a3)<=(!b5))));
  assign y12 = (((3'sd2)*(p6?p5:p5))?(3'd1):((4'd3)?(b1^~p12):(b5!==a3)));
  assign y13 = (a2!==b4);
  assign y14 = $signed(((p0>=p13)<<(p17-p11)));
  assign y15 = (((|(~a1))<<<(a4^~a4))?((2'd2)?(-5'sd3):(^p8)):((a2?b2:a1)?(~b5):(a2&a4)));
  assign y16 = $unsigned((5'd18));
  assign y17 = ((((5'd10)<<<(-(~&b1))))&(5'd27));
endmodule
