module expression_00517(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({{(5'd19),(4'd3),(4'd2)}}?{((4'd7)?(3'd4):(4'sd0))}:((-5'sd12)!=(3'sd3)));
  localparam [4:0] p1 = {(-4'sd0),(-5'sd9),(5'd21)};
  localparam [5:0] p2 = {(2'd3),{(-3'sd2)},((-4'sd6)>>>(5'd15))};
  localparam signed [3:0] p3 = (((-5'sd10)?(-2'sd0):(-3'sd1))>=(2'd1));
  localparam signed [4:0] p4 = ((((4'd12)^(5'd13))?((2'sd1)>=(5'sd11)):(!(5'd23)))<<<({2{(3'd1)}}?((4'sd0)>>>(-5'sd12)):((5'sd13)!=(4'd1))));
  localparam signed [5:0] p5 = (&(+((2'd1)==(-4'sd7))));
  localparam [3:0] p6 = ({1{(((5'd16)!==(2'sd0))||((4'sd4)!=(5'd5)))}}|((4'd1)<<((2'd3)>(5'sd7))));
  localparam [4:0] p7 = (+(^(~|(&(~|(2'd1))))));
  localparam [5:0] p8 = ((5'sd3)<=(5'd24));
  localparam signed [3:0] p9 = (5'd24);
  localparam signed [4:0] p10 = {4{(5'd3)}};
  localparam signed [5:0] p11 = (-(!(5'd2 * ((4'd13)==(2'd1)))));
  localparam [3:0] p12 = {(((4'd0)?(-2'sd0):(2'd3))==(3'd6)),{(4'd15),(2'sd0),(2'd0)},(4'sd2)};
  localparam [4:0] p13 = ((2'd0)||(2'd2));
  localparam [5:0] p14 = ({1{((5'sd3)?(2'sd1):(-2'sd1))}}?{1{((2'd0)?(4'sd5):(5'd17))}}:((2'd2)&(3'd4)));
  localparam signed [3:0] p15 = {2{(((5'd17)?(2'd3):(3'd4))?((5'sd1)?(5'd31):(3'd7)):{2{(5'd31)}})}};
  localparam signed [4:0] p16 = (6'd2 * ((5'd22)^~(2'd3)));
  localparam signed [5:0] p17 = {(3'd0)};

  assign y0 = ((~(~(&(-3'sd1)))));
  assign y1 = (((^a1)?(a5?b5:b2):(3'sd3))?(~&(4'd0)):(4'd1));
  assign y2 = (-$unsigned({4{(|(a0==b3))}}));
  assign y3 = {4{{4{p2}}}};
  assign y4 = {(!(b4?p6:a5)),(+{{a3,p5}}),(b0?a5:a1)};
  assign y5 = ({p9,p2}?(2'd2):{p14,p5});
  assign y6 = ((~^a2)?(3'd7):(a3));
  assign y7 = $signed((^(|(~|(($signed((~|b3))?{p16,a1}:(&(b2?a2:p15))))))));
  assign y8 = {({p2,p9,b3}?(p17?b4:p12):(a4?b3:p9)),{(a0?p15:b2),(p10?b3:p16)}};
  assign y9 = (3'd1);
  assign y10 = (((&(-2'sd1))>>(p14%p16))==($signed((~|p10))&(~(~p2))));
  assign y11 = {((!b5)===(a0^~a2)),{{1{p17}},(b5||p0)}};
  assign y12 = (p13<<<p11);
  assign y13 = (+{(-$signed((~|{(6'd2 * (~&p14)),(~^(a0^~p12))})))});
  assign y14 = (!((&b5)?(|p1):(b5?a3:p9)));
  assign y15 = {3{{3{b2}}}};
  assign y16 = ({$unsigned({b4,b1})}<<<((a0+b4)||(b4>>>b0)));
  assign y17 = {$signed($unsigned($unsigned(((-3'sd2))))),(-(5'd2 * (b2===a0))),{1{$unsigned({1{(~{p16,p4})}})}}};
endmodule
