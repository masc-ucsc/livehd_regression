module expression_00760(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(^(~(+(!(!(^(~|(|(-(|(|(&(|(4'd8)))))))))))))));
  localparam [4:0] p1 = (^(-3'sd0));
  localparam [5:0] p2 = (4'sd3);
  localparam signed [3:0] p3 = ((-5'sd12)-((~&(4'd11))+((5'sd13)!==(2'd0))));
  localparam signed [4:0] p4 = {4{((3'd4)?(2'sd0):(2'sd1))}};
  localparam signed [5:0] p5 = (^(&{{(~(-3'sd2)),(^(-4'sd3))}}));
  localparam [3:0] p6 = (-(((2'd0)|(2'sd1))&&(^(-3'sd3))));
  localparam [4:0] p7 = ((3'd5)===(5'd27));
  localparam [5:0] p8 = {(-{(5'd14),(4'd12),(5'd28)}),(!((2'd1)>=(5'd9)))};
  localparam signed [3:0] p9 = ({4{(3'd2)}}^~((5'sd12)>>((-3'sd2)?(2'sd1):(-4'sd2))));
  localparam signed [4:0] p10 = ((~^(((-4'sd3)?(-2'sd1):(5'd29))^(5'd2 * (5'd27))))?(((2'd2)^~(4'd2))!==(5'd14)):(~(~(!(4'd11)))));
  localparam signed [5:0] p11 = ((-((|(3'd1))<(~|(5'd26))))^(|(~|((~|(3'd5))&((5'd25)&(2'sd0))))));
  localparam [3:0] p12 = ((4'd0)<<(^(-4'sd4)));
  localparam [4:0] p13 = (((5'd15)*(-4'sd3))>>((4'd5)>>>(-3'sd3)));
  localparam [5:0] p14 = (-((((2'd0)-(-3'sd0))&&(+(4'd6)))^((5'd9)?(2'sd0):(3'd1))));
  localparam signed [3:0] p15 = (&(~{((2'sd0)?(-3'sd3):(5'sd2)),{{(3'd7),(5'd22)},{(3'd5),(5'sd11),(2'd2)}},{(-3'sd3),(3'd0),(2'd3)}}));
  localparam signed [4:0] p16 = ({2{(-2'sd0)}}|{2{(3'd5)}});
  localparam signed [5:0] p17 = {4{(-3'sd3)}};

  assign y0 = ((4'sd7)+((p13%p3)/p17));
  assign y1 = (|({(b0===b3),{3{b0}},(~|a1)}>=(~&((b1>=b3)^~(b5-p17)))));
  assign y2 = $signed(({p8,p8,p0}));
  assign y3 = {p13,p3,p12};
  assign y4 = (((b2?b2:a4)!==(~&a3))<<{4{p7}});
  assign y5 = ((+(~&b4))>>(!(+a5)));
  assign y6 = (~^(3'sd1));
  assign y7 = ((3'sd0)>=(5'd7));
  assign y8 = (5'd2 * a2);
  assign y9 = $signed(((a4%b0)/p0));
  assign y10 = (5'd2 * {1{(^a0)}});
  assign y11 = ((5'd21)?({b1,p7,a2}?(b4||a2):(2'sd1)):(5'sd13));
  assign y12 = (b2?a3:a4);
  assign y13 = $signed((5'd6));
  assign y14 = (!(|$unsigned(p13)));
  assign y15 = (((+b1)?(p0>=a5):(a1>=b4))||(-(~|((~|b5)>=(-b4)))));
  assign y16 = $unsigned($signed((((+p15)&$unsigned(p16))<=(+(a5==p0)))));
  assign y17 = ((~|(((b3?a2:a4))?($signed(a3)):(b4^~b1))));
endmodule
