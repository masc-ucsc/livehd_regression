module expression_00295(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({{3{(2'sd1)}},{(-4'sd4)}}|(((4'd12)>>>(5'd19))&{4{(3'd3)}}));
  localparam [4:0] p1 = {4{{(2'sd0),(5'd20),(2'sd1)}}};
  localparam [5:0] p2 = (((3'sd0)?(-4'sd4):(3'sd0))?{1{(5'd20)}}:{1{(4'd3)}});
  localparam signed [3:0] p3 = (5'd8);
  localparam signed [4:0] p4 = {1{((^(-4'sd5))==(|(4'sd7)))}};
  localparam signed [5:0] p5 = (-5'sd9);
  localparam [3:0] p6 = (((-4'sd6)|(2'sd0))-(|(4'd12)));
  localparam [4:0] p7 = ((2'd1)===(5'd8));
  localparam [5:0] p8 = (-3'sd1);
  localparam signed [3:0] p9 = (4'd2 * ((4'd2)<<(5'd1)));
  localparam signed [4:0] p10 = ((3'sd2)?(5'd27):((-4'sd0)?(-4'sd7):(4'd9)));
  localparam signed [5:0] p11 = (|(((+(-5'sd15))+(~&(5'sd0)))===((4'sd7)?(2'd0):(3'd6))));
  localparam [3:0] p12 = (-5'sd2);
  localparam [4:0] p13 = ((((3'd4)-(-4'sd7))|((4'd10)<=(4'sd2)))>(((3'sd2)<=(5'd5))<=((-2'sd0)<<(4'sd1))));
  localparam [5:0] p14 = {({1{{1{(2'd3)}}}}^(~|((3'd2)!==(4'sd1))))};
  localparam signed [3:0] p15 = {(3'sd0),(4'd1)};
  localparam signed [4:0] p16 = ((+(^(+(4'd14))))|(~|(|((5'sd7)?(4'd5):(5'd18)))));
  localparam signed [5:0] p17 = (^(~&{(2'd1),(3'd3)}));

  assign y0 = ((((p10?p0:p10)?(b2?p4:p7):(p6?b0:p14)))&&({p7,b3}?(a1|a2):(a5<<p17)));
  assign y1 = ((~(4'd4))-({b1,a1}==(+a5)));
  assign y2 = (~&b3);
  assign y3 = $signed((|((-2'sd1)?(-4'sd4):(b4?p14:p0))));
  assign y4 = ((3'd6)?({a4,b2}+(b1!==b0)):{4{(a1|a0)}});
  assign y5 = $unsigned((2'sd1));
  assign y6 = {b2,p11};
  assign y7 = (a3|p11);
  assign y8 = (&((b5||a3)^~{b0,b0}));
  assign y9 = (-({{(p12^p11)},{(p10>>p0)}}+(~{3{{{3{p14}}}}})));
  assign y10 = (p8||a5);
  assign y11 = (((a5-b1)!={p6,a3,p14})^(!{(p17==p16)}));
  assign y12 = {4{{1{p2}}}};
  assign y13 = (&(|((p15>>p6)?(a5!=b1):(a0?b5:p16))));
  assign y14 = (5'd28);
  assign y15 = {$signed((((+{p4,p1})&&(^(^(p2?p6:p6))))))};
  assign y16 = (~|(&(&$unsigned(((p2-p9)||$unsigned(p3))))));
  assign y17 = {3{{4{p16}}}};
endmodule
