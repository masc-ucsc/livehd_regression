module expression_00281(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-(+(|{1{(~(5'd9))}})))|({4{(3'd2)}}>((5'd20)||(5'd7))));
  localparam [4:0] p1 = (((~^((5'd30)>(4'd9)))<((-3'sd1)>=(-2'sd1)))!==(~&(3'd1)));
  localparam [5:0] p2 = (!((&(-4'sd6))?(~|((-5'sd14)|(4'sd4))):(-(-2'sd1))));
  localparam signed [3:0] p3 = {3{((^(2'd3))&&{2{(2'd2)}})}};
  localparam signed [4:0] p4 = (-(6'd2 * (5'd2 * (5'd17))));
  localparam signed [5:0] p5 = ((-4'sd5)?((4'd1)<<(2'd2)):{(3'd5),(-4'sd2)});
  localparam [3:0] p6 = (4'd2 * ((3'd1)^(4'd7)));
  localparam [4:0] p7 = (3'sd2);
  localparam [5:0] p8 = (((5'd22)^(2'd0))?((3'd2)|(3'd4)):((4'd6)<<<(-3'sd1)));
  localparam signed [3:0] p9 = ({1{{(3'd1)}}}!==((-5'sd14)+(5'd3)));
  localparam signed [4:0] p10 = ((6'd2 * (~|(!(5'd11))))==(~|(((5'd19)==(2'd0))<<<((-3'sd3)!==(-2'sd1)))));
  localparam signed [5:0] p11 = {2{(&(4'sd5))}};
  localparam [3:0] p12 = {(3'd7),(2'sd0)};
  localparam [4:0] p13 = {(~&{(-(+(-2'sd0)))}),{{(-2'sd1),(2'd2),(5'd25)},{(3'd4),(-4'sd3)}},(^{{(-2'sd0),(4'd10)},(&(4'd12))})};
  localparam [5:0] p14 = (+(!(~|((&(5'sd15))||(~(-2'sd1))))));
  localparam signed [3:0] p15 = (((5'd7)>(3'd0))%(4'd6));
  localparam signed [4:0] p16 = (3'd6);
  localparam signed [5:0] p17 = ((5'd12)!==(3'd7));

  assign y0 = (&(a4?a5:a2));
  assign y1 = (({4{p9}}==(&(a4<<<p17)))|(|((p7<<p2)?(~&{3{b4}}):(p1?p13:b0))));
  assign y2 = {4{{4{b3}}}};
  assign y3 = {1{({({3{b3}}),(4'd5)}!=$signed((~&({4{a5}}==(b5==b1)))))}};
  assign y4 = (~&(~&((~(!(~&p16)))>>>(~|(^(p7*p2))))));
  assign y5 = {({1{{($unsigned(p8)),{2{p17}}}}}==(-{2{((^a2))}}))};
  assign y6 = ({3{{b0,p5}}}|{3{{a5}}});
  assign y7 = (({4{p1}}||(p8?p11:p10))|((p16^p13)<<<(p2?p10:b5)));
  assign y8 = {((-4'sd5)!=(3'd2)),({p15,p6}<<(p11>p12)),(5'd5)};
  assign y9 = (((3'd3)?(b4^~b1):(~^(3'd7)))>((5'd21)>(|(4'd0))));
  assign y10 = ({{(p8>>>b5),(a0===b1),(p14&p0)}}<<((6'd2 * a2)>>>(4'sd1)));
  assign y11 = (a0&b1);
  assign y12 = (((p6!=p12)||(p11?b0:a1))?((a1!=a1)||(a0?p6:p14)):{(a3?a0:b1),{2{b3}}});
  assign y13 = (($unsigned((~(3'd0))))<<((5'd2 * p7)?(!(a1||b5)):(p3==p11)));
  assign y14 = {$unsigned($unsigned(p7))};
  assign y15 = ((~|(!(-2'sd1)))<<<((~|p2)?(-5'sd14):(4'd13)));
  assign y16 = {({((a3?b1:b0)===(b2&a4))}?{2{{4{a5}}}}:((a3&b4)?{b4,p3,a0}:{1{b4}}))};
  assign y17 = (!$unsigned((~|(|(5'd12)))));
endmodule
