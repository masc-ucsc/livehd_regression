module expression_00473(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'd2)?(-4'sd6):(4'd15))|((4'd0)<(-4'sd2)));
  localparam [4:0] p1 = ((4'd12)?(-2'sd0):((3'd3)?(2'sd1):(3'd2)));
  localparam [5:0] p2 = ((|((^(-(3'sd0)))<<<((2'd3)>(4'sd2))))+(((-2'sd0)*(4'd3))>((3'sd3)<=(-4'sd5))));
  localparam signed [3:0] p3 = (3'd6);
  localparam signed [4:0] p4 = (4'd2);
  localparam signed [5:0] p5 = (!(^(~|(~^(~|(!(+(~(^(~^(-(-(&(-3'sd1))))))))))))));
  localparam [3:0] p6 = ((((5'sd10)<<<(-4'sd7))>>((-2'sd1)<(-4'sd4)))+((-(5'd2))!=((3'd2)==(-5'sd0))));
  localparam [4:0] p7 = {2{(2'd1)}};
  localparam [5:0] p8 = (-4'sd1);
  localparam signed [3:0] p9 = (((5'sd7)?(3'd5):(3'd5))^((2'sd1)>>>(3'sd2)));
  localparam signed [4:0] p10 = (((4'd6)!==(2'sd1))|{3{(2'd3)}});
  localparam signed [5:0] p11 = (!(~^((|(~^((-5'sd12)^~(3'd3))))||(!(!(~^(2'd3)))))));
  localparam [3:0] p12 = ((((3'd4)||(2'd2))^~((3'd2)/(5'sd2)))>>(((-5'sd13)?(2'd0):(-3'sd3))!=((-4'sd3)|(5'd8))));
  localparam [4:0] p13 = (~^(6'd2 * {(5'd8),(4'd13),(5'd0)}));
  localparam [5:0] p14 = ((~^((~|(-(5'd4)))&&{4{(2'sd0)}}))+{1{(-2'sd1)}});
  localparam signed [3:0] p15 = ((~|(!((-3'sd0)?(-4'sd0):(-5'sd15))))?(6'd2 * (|(2'd0))):(((5'd21)!=(2'd1))!={(2'd3),(2'sd0),(3'd5)}));
  localparam signed [4:0] p16 = ((3'd4)!=({4{(-2'sd0)}}==={3{(2'sd0)}}));
  localparam signed [5:0] p17 = {1{{3{((5'd8)?(5'd0):(3'd4))}}}};

  assign y0 = {(~&({(p1^p17),(p10>>>p10),{p0,p17,a5}}?({p0,p15,p9}>=(4'd3)):{(~^p16),(-p15),(p11?p0:p6)}))};
  assign y1 = (((6'd2 * p13)<<{p10,p7,p2})<<(4'd15));
  assign y2 = ($signed(((b2<<a2)>(b3==b0))));
  assign y3 = {((b3)?(a4+b0):{p12,p9,p16}),(-4'sd7),((b3>>p15)>>>(a2<a5))};
  assign y4 = (~|b0);
  assign y5 = ($signed(((~&((^p17)?(~^p4):(^p10)))?(|(|$unsigned((p13?p9:p12)))):(|{3{{4{p9}}}}))));
  assign y6 = (2'd2);
  assign y7 = (!(-(5'd25)));
  assign y8 = (({$unsigned(p10)})?((b1?a0:p4)):((a2+a5)!==(b3===b1)));
  assign y9 = ((((&b3)!==(a2^b3))<(|(b5?a2:a4)))<((^(b2+b2))*(^(a4<=a1))));
  assign y10 = ($unsigned((^{{b1},(5'd2 * a0)}))<<<(^{$unsigned({b3,b2})}));
  assign y11 = ((-4'sd6)<={(b5?p5:p14)});
  assign y12 = (5'sd10);
  assign y13 = ((+b1)&&(a1));
  assign y14 = {((p7<<p7)<<<(b5&a3)),(5'd2 * (b1?a2:b0))};
  assign y15 = (&((&((b1?p7:a1)^~(a3?b0:b2)))?(+(~&(-2'sd0))):((+a1)?(2'd1):(p12>=b1))));
  assign y16 = {(b1^~p8),{2{a1}}};
  assign y17 = (~$signed($unsigned({4{(4'd12)}})));
endmodule
