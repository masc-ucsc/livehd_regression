module expression_00573(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd19)^~(-3'sd2));
  localparam [4:0] p1 = (|(((~^((5'd28)<<(4'sd7)))+(~|(&(4'd10))))>=((&((3'd6)-(-4'sd0)))>>(&(&(5'd17))))));
  localparam [5:0] p2 = (~|{{(~{(4'sd0),(5'd10)})},(~^(^{(5'd19)})),(|(~&(^(-3'sd2))))});
  localparam signed [3:0] p3 = (~{(5'sd10)});
  localparam signed [4:0] p4 = (({(2'sd0),(5'd29),(4'd12)}>(((2'd1)?(-4'sd2):(5'sd7))||{(2'd2)}))>={((2'd2)?(-5'sd5):(3'sd0)),((4'd3)?(3'd4):(3'd2)),{((-2'sd1)>>(5'd10))}});
  localparam signed [5:0] p5 = (&((2'sd0)<(4'd3)));
  localparam [3:0] p6 = {((-4'sd7)?(3'd6):(4'd8)),((4'sd2)?(2'sd1):(2'sd0)),{1{(4'd6)}}};
  localparam [4:0] p7 = ((4'sd1)-((3'd2)<=((5'd31)+(-(-3'sd1)))));
  localparam [5:0] p8 = {{3{({(3'sd3)}==((-5'sd5)==(5'd12)))}}};
  localparam signed [3:0] p9 = {2{{4{(2'sd1)}}}};
  localparam signed [4:0] p10 = ((3'd1)<=(3'd4));
  localparam signed [5:0] p11 = ((-2'sd1)>>(2'd3));
  localparam [3:0] p12 = ((((5'sd5)<<<(3'sd0))&&{(2'd2),(3'sd1),(-2'sd1)})>({(-3'sd1),(4'd15),(4'sd0)}<<((2'd2)<(3'd4))));
  localparam [4:0] p13 = ((+(((-5'sd4)|(-3'sd2))-((4'd4)>>(3'sd2))))!=(((4'd15)?(5'd29):(2'sd0))?((-2'sd1)%(2'd0)):(^((3'd6)?(4'd11):(2'd1)))));
  localparam [5:0] p14 = (~|((~{1{(-2'sd0)}})==((5'd11)?(-4'sd5):(5'd4))));
  localparam signed [3:0] p15 = {4{((-2'sd0)?(5'd0):(-2'sd0))}};
  localparam signed [4:0] p16 = {{{(2'd3),(-2'sd0)},((-5'sd0)^~(4'sd6))},{(2'sd1)}};
  localparam signed [5:0] p17 = (&(+((4'd13)&&(3'd2))));

  assign y0 = (b2?p14:p3);
  assign y1 = ((b2?b1:p9)?{b5,b2}:(3'd5));
  assign y2 = $signed($signed((b3?p11:a1)));
  assign y3 = ({b0}?(p3!=b0):{3{p16}});
  assign y4 = ($signed((+((-(+(!p12)))>>>(^(~$signed(p3))))))>=(+((~|(|(a0&a2)))<<<((a3)+(&p14)))));
  assign y5 = (((a2===b0)<<(a4*b2))!=($unsigned(a0)?$signed(a3):$signed(b3)));
  assign y6 = ((3'sd3)&&(5'd14));
  assign y7 = ({a2,b0}+(b4==b4));
  assign y8 = (5'd26);
  assign y9 = (4'd3);
  assign y10 = {4{p7}};
  assign y11 = $signed($unsigned(a3));
  assign y12 = {2{{3{$signed((a0^~a2))}}}};
  assign y13 = (-5'sd0);
  assign y14 = {{{2{p0}}},{{p3},(|p10)},{2{(|p12)}}};
  assign y15 = ((p16?b3:p3)+(-2'sd1));
  assign y16 = ((((~&b1)||(b5+b2))&({b1,b1}>>$unsigned(a0)))!==((~(4'd2 * (~&$unsigned(a4))))));
  assign y17 = ((((a3<<a1)===$signed(a0))==({1{p5}}>(-a4)))>={2{(~&(-(a4<<b1)))}});
endmodule
