module expression_00424(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd2);
  localparam [4:0] p1 = ((~{1{({3{(-2'sd0)}}+((3'd0)<<(5'sd12)))}})=={1{(((4'd7)<<(-3'sd3))=={3{(3'sd1)}})}});
  localparam [5:0] p2 = (((3'sd2)?(-2'sd1):(4'd2))?((4'd4)?(5'd7):(5'd18)):(((5'sd11)>=(3'sd3))&&((4'd12)?(3'd1):(4'd9))));
  localparam signed [3:0] p3 = (((4'sd1)?(4'd0):(-4'sd0))?((3'd0)^(-2'sd0)):((4'd5)?(-3'sd1):(4'sd2)));
  localparam signed [4:0] p4 = {((-3'sd1)>(-2'sd0)),((5'd23)?(5'd14):(3'sd1)),{(-3'sd2),(4'sd3),(-4'sd7)}};
  localparam signed [5:0] p5 = (~&((3'd2)!==(4'd4)));
  localparam [3:0] p6 = ({2{((2'sd0)||(4'sd7))}}<=(2'd1));
  localparam [4:0] p7 = (-2'sd1);
  localparam [5:0] p8 = (-((-5'sd5)!==(-((4'sd7)==(^(2'sd0))))));
  localparam signed [3:0] p9 = {4{((4'd11)<(2'sd0))}};
  localparam signed [4:0] p10 = (^((3'd2)!=(4'd7)));
  localparam signed [5:0] p11 = ((5'd16)?(4'sd3):((4'd4)?(-3'sd2):(5'sd10)));
  localparam [3:0] p12 = (~({4{((4'sd2)?(5'd20):(2'sd0))}}>({4{(-4'sd0)}}>>(&{1{(5'd11)}}))));
  localparam [4:0] p13 = (!((&(+(3'sd2)))?((2'sd1)>>(4'd2)):(+(~&(-5'sd5)))));
  localparam [5:0] p14 = (!(~&((~|(5'd13))&&(~|(4'sd4)))));
  localparam signed [3:0] p15 = ((5'd6)?(5'd18):(-5'sd13));
  localparam signed [4:0] p16 = ((((-5'sd7)==(4'd9))&((2'd2)<(3'd5)))||({(-3'sd0),(5'd31),(5'd6)}-((-3'sd3)<<<(-3'sd3))));
  localparam signed [5:0] p17 = ((4'd2 * ((3'd7)+(3'd4)))>>>(6'd2 * ((5'd4)!==(3'd5))));

  assign y0 = (-3'sd2);
  assign y1 = ((2'sd0)<(2'd2));
  assign y2 = {({4{(b4==b1)}}<={1{({a0,a2}<<<(a2-b5))}})};
  assign y3 = {(2'd2)};
  assign y4 = (5'd3);
  assign y5 = ((p12==p0)?(b4<=p0):(p8?p6:a5));
  assign y6 = (3'd1);
  assign y7 = {(3'sd3),{a4,p6,p0}};
  assign y8 = {((3'd0)?(5'd17):(b2>p7))};
  assign y9 = {1{{3{{4{p10}}}}}};
  assign y10 = (&((5'd14)>>>((3'd4)!={2{(2'sd0)}})));
  assign y11 = (p8^b0);
  assign y12 = (-((3'd2)&$unsigned((~|(-2'sd0)))));
  assign y13 = {1{(2'sd0)}};
  assign y14 = {1{{1{(p2^a0)}}}};
  assign y15 = ((p10<<a5)-(!(b4&&p16)));
  assign y16 = (-3'sd0);
  assign y17 = (~|(((|(^(~^a5)))<<<(4'd2 * (~^b0)))>={1{{3{(a5!==a2)}}}}));
endmodule
