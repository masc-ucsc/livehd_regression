module expression_00220(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{3{{1{((4'd13)&(2'sd0))}}}}};
  localparam [4:0] p1 = {1{{{((2'd1)?(4'sd5):(4'sd3)),((3'd1)?(4'd5):(5'sd13)),{(-2'sd1),(4'sd7)}}}}};
  localparam [5:0] p2 = ((3'sd1)%(3'sd0));
  localparam signed [3:0] p3 = ({3{(3'd7)}}==(((2'd3)+(5'd2))>=((2'sd1)>>(2'sd0))));
  localparam signed [4:0] p4 = (&(&(-3'sd0)));
  localparam signed [5:0] p5 = ((((~&(2'd2))^{1{(-5'sd3)}})-(6'd2 * {3{(5'd19)}}))||{2{(((-5'sd6)==(3'd1))<<<((5'd3)!=(5'd16)))}});
  localparam [3:0] p6 = {{(^{3{(5'd13)}}),(~&{(3'sd3)})},{{(-5'sd3),(4'd7),(3'd7)},{4{(5'sd5)}}}};
  localparam [4:0] p7 = (~&(((~&(2'sd1))?((2'd2)^~(4'd14)):((-3'sd1)^~(4'd12)))===(((5'd25)?(3'd1):(-5'sd7))?((3'sd1)?(2'd2):(5'd4)):((-4'sd1)?(-5'sd5):(5'sd10)))));
  localparam [5:0] p8 = {((((4'd15)>=(2'sd0))-{(4'sd4),(4'd7)})^~(((5'sd7)>>(5'sd13))<={(4'd10),(4'd14)}))};
  localparam signed [3:0] p9 = (~{2{(~|{4{(-2'sd1)}})}});
  localparam signed [4:0] p10 = ((5'd28)===(5'sd10));
  localparam signed [5:0] p11 = (~^{3{((+(-3'sd0))==(~|(2'sd0)))}});
  localparam [3:0] p12 = (&(((2'sd1)<<<(-4'sd7))>=((5'd11)+(5'd14))));
  localparam [4:0] p13 = {1{{2{{4{(3'd2)}}}}}};
  localparam [5:0] p14 = {(~|(^{(-2'sd0),(2'd2),(5'd14)})),{{(4'sd4),(5'd11)},{(3'sd0),(5'sd10),(2'd1)}},{(&{(3'd1),(5'd26),(-4'sd3)})}};
  localparam signed [3:0] p15 = (5'd15);
  localparam signed [4:0] p16 = (4'd14);
  localparam signed [5:0] p17 = ({((3'd2)?(-2'sd1):(-4'sd7))}?(-2'sd0):((4'd10)?(-4'sd0):(-4'sd4)));

  assign y0 = ((p1?a4:a2)%a0);
  assign y1 = {(~^(-{p13,p10})),{(~&p11),(!p1)},{p1,p14,p7}};
  assign y2 = {1{(^$signed({2{$signed(($signed(($unsigned({4{p14}})))))}}))}};
  assign y3 = (p15?p5:a2);
  assign y4 = (!(^{{p4,a0},(~&$unsigned(p17))}));
  assign y5 = (4'd13);
  assign y6 = (!(3'sd0));
  assign y7 = (4'd1);
  assign y8 = {2{(-(p8+a1))}};
  assign y9 = {({(a3>=a0)}<<<{p13,b0,p9}),{((a5^p7)>{b0})}};
  assign y10 = (4'd2);
  assign y11 = (~&((((-(~&b1)))!=(^(!(+p13))))<=(3'sd0)));
  assign y12 = {{(~|p2),(+p11),{a4,a3,a0}}};
  assign y13 = {(&(^(({p8,p11}>={a0,p15,p9})-{((p0?p11:p10)?(p7>p12):(p3<=p5))})))};
  assign y14 = ({(p2?b1:a2),(a3?a3:a3),{a2,a4,p13}}?{{a0,a4},(a4?a2:b0)}:((a0<<<p10)?(b1?a0:b3):{b0,a0,p7}));
  assign y15 = (((~&(5'd2 * (5'd8)))>=$unsigned((~^(^(a2^~b1)))))||((5'd9)!=((3'd6)==(p14!=p4))));
  assign y16 = (|(+(!{(~&{(~&(-p1)),{p16,p14}}),{(|b4),{p5},(~^p14)}})));
  assign y17 = $signed(a2);
endmodule
