module expression_00586(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{{2{((5'sd11)+(3'sd2))}}}}?({(-2'sd0)}?(|(5'd1)):(~&(5'sd10))):((-(5'd11))?((2'd0)<<<(2'd1)):((4'd15)-(2'sd1))));
  localparam [4:0] p1 = {{(2'd2),(-2'sd0),(-4'sd7)},{{1{((4'sd2)>>>(2'sd1))}}},{4{(2'sd0)}}};
  localparam [5:0] p2 = (2'sd1);
  localparam signed [3:0] p3 = {{((3'd7)<<(4'd12)),((5'd20)>=(-5'sd5)),{(2'd3)}}};
  localparam signed [4:0] p4 = (3'sd0);
  localparam signed [5:0] p5 = (+(5'd26));
  localparam [3:0] p6 = (((4'sd2)?(-2'sd1):(3'sd0))?((5'd25)?(3'sd1):(4'd10)):((5'd30)?(5'd25):(-2'sd1)));
  localparam [4:0] p7 = (!(5'd22));
  localparam [5:0] p8 = (-({{(4'd0),(4'd2),(3'sd3)}}&&(^{(2'd1),(4'd9),(5'sd14)})));
  localparam signed [3:0] p9 = {({((5'd12)^~(-3'sd2)),((4'd14)?(3'd3):(3'sd1))}?{(~|(-3'sd2)),(-(5'd2))}:((3'd0)?(-5'sd5):(3'd7)))};
  localparam signed [4:0] p10 = {{2{({4{(5'd13)}}<={3{(4'sd0)}})}}};
  localparam signed [5:0] p11 = (~^(5'd2 * (2'd3)));
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = {4{{1{(&(2'd3))}}}};
  localparam [5:0] p14 = {3{(~((2'd3)||(2'd1)))}};
  localparam signed [3:0] p15 = (~^{1{(5'd20)}});
  localparam signed [4:0] p16 = ((+{1{(~(2'sd0))}})!=(((2'd2)<(2'd1))&&((5'd13)|(-3'sd0))));
  localparam signed [5:0] p17 = (2'sd0);

  assign y0 = {{(b3!==b5),(p7?a2:p10),(5'd2 * p8)}};
  assign y1 = (3'd5);
  assign y2 = (2'sd1);
  assign y3 = ((3'sd2)-(~|(2'd2)));
  assign y4 = ((((a4!==a1)===$unsigned(a0))>>>(((b1==p14)|$signed(b2)))));
  assign y5 = (((p0>a3)-{1{(-4'sd4)}})>((p11>p4)+(a3&&b4)));
  assign y6 = {(a4>>p15)};
  assign y7 = (~{a2,b5});
  assign y8 = {2{(4'sd0)}};
  assign y9 = (((p0&&a3)?(~^p15):(a3/p11))^((-5'sd6)*(p6+a2)));
  assign y10 = $unsigned((4'd11));
  assign y11 = {{2{(-p0)}},{{4{b0}}},({2{p6}}<<{2{b0}})};
  assign y12 = (~^$unsigned(((^{(&{b4,b2,b4}),({b2}<<(-b2))})|$unsigned((4'd2 * $unsigned((~b5)))))));
  assign y13 = (-((!(4'd11))^(2'd3)));
  assign y14 = (((-2'sd1)^({p1,a5,a3}|$signed(a3)))!=$signed((3'sd1)));
  assign y15 = (~^(~^$signed((((a3!=b0)-(p10<<<p13))+(|((|p8)+{2{a2}}))))));
  assign y16 = ({((a1!==a0)==(b2-a0)),({a5,p9,p15}+(p13-p13))}>={((p3<<a5)!={(b3>>>p0)})});
  assign y17 = (^({{a1,a1,p17},(~|b2),(b5<<<a3)}<<<{(b2===b4),(b2^~b3),(b2>b5)}));
endmodule
