module expression_00455(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-((5'd25)?(^((5'd2)||(5'd31))):(~|(-(-2'sd1)))));
  localparam [4:0] p1 = ({(4'sd6),(2'd1),(-3'sd1)}^(3'd1));
  localparam [5:0] p2 = (({3{(2'd1)}}>(~&(3'd5)))<={((4'd13)>=(3'sd3)),{(4'd2),(3'd0),(-2'sd0)},((2'd3)?(3'd3):(3'd6))});
  localparam signed [3:0] p3 = {{3{(-5'sd5)}},(((3'd0)^(-4'sd7))!={3{(-5'sd14)}})};
  localparam signed [4:0] p4 = ({1{({{(-3'sd0)}}&&{1{{1{(-4'sd4)}}}})}}>{1{(4'd2 * {3{(3'd4)}})}});
  localparam signed [5:0] p5 = (((~|(~^(-4'sd2)))<<<(&((5'd21)-(5'sd8))))<=((&((3'd0)<<(-4'sd2)))!=((4'sd0)<=(-3'sd3))));
  localparam [3:0] p6 = {4{((5'd18)>(3'd7))}};
  localparam [4:0] p7 = (-4'sd4);
  localparam [5:0] p8 = ((-(4'sd5))==((4'd9)||(2'sd1)));
  localparam signed [3:0] p9 = (((3'd6)>>>(3'd3))?((5'd7)?(4'd13):(2'd0)):((-4'sd3)?(2'd0):(2'sd0)));
  localparam signed [4:0] p10 = (((-4'sd4)+(4'sd5))>=((4'd15)?(2'sd0):(2'd0)));
  localparam signed [5:0] p11 = (~|(((4'd11)&(-2'sd1))>>>((5'd18)<<<(3'd7))));
  localparam [3:0] p12 = (~((((4'sd1)<=(5'd15))<<((2'd2)&(4'd12)))>(+((~|{2{(3'd1)}})>(&((3'sd0)?(5'd23):(-5'sd1)))))));
  localparam [4:0] p13 = (+{(((3'sd1)>=(4'd4))?(~&(5'd23)):((3'sd3)<<<(2'd3))),(((5'd21)&&(3'd6))?((5'sd5)<<(3'sd2)):((4'd13)>>>(4'd7)))});
  localparam [5:0] p14 = (((4'sd0)?(2'd3):(2'd2))|{1{(5'd18)}});
  localparam signed [3:0] p15 = {4{(-2'sd1)}};
  localparam signed [4:0] p16 = (((5'sd4)?(3'd2):(4'd3))?(~^(~^(&(-5'sd15)))):(~^((5'sd4)?(-5'sd14):(4'd2))));
  localparam signed [5:0] p17 = (((2'd3)===(2'd0))^~(~^(~^(((2'sd0)/(-4'sd5))>(4'd8)))));

  assign y0 = ({((&{{p4,b5,p17}})>>>(5'd13))}>>>{(!(~^b2)),(b2!==a3),(3'd2)});
  assign y1 = {1{{1{$signed((~{2{p17}}))}}}};
  assign y2 = ((((p6!=a2)?(p0?a0:p3):(a4?a1:b3)))|((p15?a1:p9)&&(+(&b5))));
  assign y3 = {(|(p2==b1)),(b0&&a2),(~(p11))};
  assign y4 = (((a5<b5)?(5'd31):{p4,p16,b1})?({a2,b2,a3}?{p2}:(p11>>>a5)):{{a3},(p4^p4)});
  assign y5 = $unsigned(({(&p3),{p1,a1,p9}}));
  assign y6 = {3{((p15||a3)|(-5'sd3))}};
  assign y7 = (3'd3);
  assign y8 = (+p1);
  assign y9 = (5'd2 * (5'd28));
  assign y10 = ((~|(4'd7))>>{(p17&a5),(b1&a5)});
  assign y11 = ((((a1&&a2)!=={4{b3}})&(~&{b5,p0}))<<<(((p11<p3)>>(b3||p8))||((a2>>>b3)||(p12^p1))));
  assign y12 = {2{p14}};
  assign y13 = (b0&&a2);
  assign y14 = ({p17,p10,p17}&&{p3,b1,p6});
  assign y15 = {1{(p1^~p17)}};
  assign y16 = (!(~^(p0?p16:p9)));
  assign y17 = ((2'sd0)===((a0?a0:b0)?(-2'sd1):(a5?b4:a3)));
endmodule
