module expression_00405(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!{(3'sd3)});
  localparam [4:0] p1 = {(4'd3)};
  localparam [5:0] p2 = ((3'd1)&(5'sd9));
  localparam signed [3:0] p3 = ((5'sd10)?{(5'd3),(3'sd0)}:(3'd3));
  localparam signed [4:0] p4 = ({{(2'd3),(-3'sd1),(-4'sd7)}}?{{(2'd0),(2'sd0)},{(-2'sd0)}}:({(-5'sd1),(2'd0)}?{(-2'sd0)}:((3'sd3)?(5'sd7):(2'sd1))));
  localparam signed [5:0] p5 = {(-(&(3'd4))),(~^((3'sd1)?(5'd1):(2'd0))),(-(~&{(5'd6)}))};
  localparam [3:0] p6 = {2{((-5'sd12)===(3'sd2))}};
  localparam [4:0] p7 = (+((2'sd1)>=(-2'sd0)));
  localparam [5:0] p8 = (~&(~(+{{(|((!(~&((4'd12)>>>(5'sd14))))^~(|{(-3'sd0),(-2'sd1),(-5'sd8)})))}})));
  localparam signed [3:0] p9 = (({1{(5'd14)}}&&{(5'd2),(-4'sd1)})?{2{{1{(-2'sd1)}}}}:{4{(2'd1)}});
  localparam signed [4:0] p10 = (((2'd0)>>>(-5'sd13))+(-5'sd11));
  localparam signed [5:0] p11 = (!(~&(3'd7)));
  localparam [3:0] p12 = (^{3{{1{{1{(4'sd4)}}}}}});
  localparam [4:0] p13 = ((~|{2{{(5'sd15)}}})^((~{4{(-3'sd1)}})===((-3'sd2)>>(3'sd3))));
  localparam [5:0] p14 = ({4{(5'd2 * (4'd14))}}&&(((3'sd0)^(-3'sd0))?((3'sd1)&&(4'd14)):((-5'sd12)?(5'd29):(4'd5))));
  localparam signed [3:0] p15 = ((((-2'sd1)?(4'd13):(2'd1))||{3{(4'sd5)}})<<<{4{(2'd3)}});
  localparam signed [4:0] p16 = ((((5'd13)<<<(3'd0))!==((5'd21)<=(4'd8)))&(((3'sd2)==(-4'sd2))&&((2'd3)-(5'sd5))));
  localparam signed [5:0] p17 = ((4'sd7)==(2'd3));

  assign y0 = (4'd0);
  assign y1 = $unsigned((-(^(4'd13))));
  assign y2 = $unsigned((($unsigned((((p16|b2))^~(p7>>>p6)))<<{2{{2{b0}}}})));
  assign y3 = $signed(((~(~$unsigned($signed((b0^~p2)))))?((+(p12?a5:p10))|$unsigned((^p5))):$signed($signed(((&b1)?(!b5):(&a0))))));
  assign y4 = (~&(4'd11));
  assign y5 = {3{(p13<<<p10)}};
  assign y6 = (!((5'sd8)?((a0?b0:p17)<(b3?b3:a3)):{a4,b1,a2}));
  assign y7 = ({1{a5}}?(p15<=p13):(a5?b4:p6));
  assign y8 = ({1{(a2?a5:a2)}}!==(-4'sd7));
  assign y9 = {((~{{1{p11}},{p11,p9,p1},{a2}})<={({p10,p4,p11}<=(p3>p2))})};
  assign y10 = (4'd10);
  assign y11 = ((((~|a1)>=(a3-b1))^~(&$unsigned((a2+b2))))!==$signed((!(((a3<<a4)-(&b4))>$unsigned((!(+b2)))))));
  assign y12 = (a4===a3);
  assign y13 = {2{p12}};
  assign y14 = (~^((p14^p13)*(p14/p15)));
  assign y15 = {(-{(|(~{1{{a4,a2,b3}}})),{3{(~&a1)}}})};
  assign y16 = (-3'sd1);
  assign y17 = (!(4'd13));
endmodule
