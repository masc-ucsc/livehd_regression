module expression_00261(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd2)?((5'd0)<<(-4'sd1)):((5'd25)?(-4'sd7):(2'd3)));
  localparam [4:0] p1 = (-5'sd15);
  localparam [5:0] p2 = {1{((((-2'sd1)?(-2'sd1):(5'd18))===((2'd3)?(3'sd3):(-5'sd12)))?(((-2'sd1)-(-4'sd6))?((5'd4)?(4'd5):(2'sd1)):{4{(3'd2)}}):(((2'sd1)?(5'sd5):(-2'sd1))?{4{(4'd13)}}:(4'd2 * (3'd4))))}};
  localparam signed [3:0] p3 = (~|(+{4{{2{(5'd11)}}}}));
  localparam signed [4:0] p4 = {{((4'sd4)>=(-3'sd1)),((3'd5)>>>(5'd19)),((-5'sd9)^~(-2'sd1))},{(|(5'sd3)),((4'sd1)?(-3'sd1):(3'sd0))},(+(!((-4'sd4)!==(4'd0))))};
  localparam signed [5:0] p5 = {3{{4{(-5'sd5)}}}};
  localparam [3:0] p6 = ((-5'sd2)?(3'sd3):(5'd24));
  localparam [4:0] p7 = ({2{(~&(~&(2'd2)))}}>(~|(&(~^(~^((-2'sd1)-(5'd12)))))));
  localparam [5:0] p8 = (~((3'd7)?(2'd1):(^((5'd5)!==(2'd1)))));
  localparam signed [3:0] p9 = ((((4'd7)?(3'sd1):(4'd13))<<((2'd1)?(4'd5):(-3'sd1)))&&{1{(((2'sd1)?(4'd12):(3'd3))?((5'sd5)-(-5'sd4)):{4{(-2'sd0)}})}});
  localparam signed [4:0] p10 = ({(3'd2),(5'sd15),(5'sd10)}||((-3'sd0)|(5'd14)));
  localparam signed [5:0] p11 = (6'd2 * ((5'd28)&(2'd2)));
  localparam [3:0] p12 = (((5'd3)+(3'd2))/(3'd6));
  localparam [4:0] p13 = {(5'sd2),{(3'd2)}};
  localparam [5:0] p14 = (!(|((&(&(((3'd5)<<(5'd14))|(-(5'd31)))))|(+(!((&(3'sd2))*(~^(3'd7))))))));
  localparam signed [3:0] p15 = (+((^(|((5'sd5)&(-4'sd6))))<<(~&(((5'd16)<<<(5'sd5))/(-4'sd3)))));
  localparam signed [4:0] p16 = (!{{{2{(4'd1)}},{(2'd0)}},(-(~^{(5'd3)})),{{(4'sd3),(5'd30)}}});
  localparam signed [5:0] p17 = ((-5'sd6)?(-3'sd2):(2'sd1));

  assign y0 = (~&(+(5'd1)));
  assign y1 = (2'sd1);
  assign y2 = (-3'sd0);
  assign y3 = (b2?p1:a1);
  assign y4 = ({2{(a5||p6)}}&({2{p10}}<(p16-b1)));
  assign y5 = (p5?p13:b3);
  assign y6 = (b1);
  assign y7 = ((&(~|p2))%p11);
  assign y8 = (p7^~p12);
  assign y9 = ((&p1)?{3{p15}}:(a2?p6:p15));
  assign y10 = $unsigned($unsigned(($signed($signed((2'd1))))));
  assign y11 = ((~^{{p10,p5},(p2<<p1),(p7&p9)})>(~(~&{(p5+p4),(&(b3>p14))})));
  assign y12 = (~^((!$unsigned((!($signed(a2)&$unsigned(p16)))))>>>(~(~^((^(-p16))>>>(a2==a2))))));
  assign y13 = {((p0?p0:p7)?(5'sd5):(p5?a0:p4)),{(-4'sd7)},(-5'sd10)};
  assign y14 = ({4{a0}}>>>((p14?p1:p16)>=(p2>p12)));
  assign y15 = ((b0<<<b1)?$unsigned({2{p16}}):(p12?p7:b2));
  assign y16 = (4'd11);
  assign y17 = (~^{((-(b0?a1:a3))?(!(a5?b3:p0)):({b1,p6,a1}?(~&b4):(-b2)))});
endmodule
