module expression_00849(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(5'sd5),(-({4{(3'd6)}}||((2'd1)&(2'sd0))))};
  localparam [4:0] p1 = {((((-2'sd0)||(-2'sd1))<=(!((5'sd15)?(2'd2):(5'sd13))))<={((4'd9)?(4'd12):(5'sd1)),((5'd27)?(2'd2):(-5'sd10)),((3'd2)?(2'd1):(3'd5))})};
  localparam [5:0] p2 = ((((2'sd1)^~(-4'sd2))^{(2'sd1),(4'd10)})>>{(~|(&(5'd8))),(~|(4'd3))});
  localparam signed [3:0] p3 = (&(3'sd3));
  localparam signed [4:0] p4 = {{{((5'd30)&&(5'd31)),(+(5'd19)),((-3'sd1)&&(5'd8))},(~^(((5'sd11)&&(-4'sd6))+((2'd1)?(5'd1):(5'd30))))}};
  localparam signed [5:0] p5 = (((((2'sd0)||(5'd12))&&((3'd0)*(2'd1)))-(((3'd3)&&(2'sd0))>=((2'd1)||(-2'sd0))))^~((((5'sd9)/(-2'sd1))%(-2'sd0))!=(((2'd2)&(3'd1))&&((4'd1)<=(3'sd0)))));
  localparam [3:0] p6 = (({(5'd27)}?(^(5'd14)):(-5'sd9))<<{3{(3'd2)}});
  localparam [4:0] p7 = (~|({4{(4'sd2)}}?(~^(-5'sd6)):((5'd14)?(5'sd9):(2'd2))));
  localparam [5:0] p8 = (~^(-5'sd2));
  localparam signed [3:0] p9 = {((2'd1)?(2'd0):(4'd0)),(~^(2'd0))};
  localparam signed [4:0] p10 = (((2'sd0)<<<(|(-5'sd10)))?(((4'd11)>(-2'sd1))!==((2'sd0)?(5'sd12):(2'sd0))):(3'd6));
  localparam signed [5:0] p11 = ({(2'd0),(-5'sd2)}?((5'sd5)<<<(2'd0)):(5'd2 * (4'd14)));
  localparam [3:0] p12 = ((2'sd0)!={((4'd2)?(5'sd2):(4'd9)),((4'sd4)>(-3'sd0)),((5'd9)|(3'd7))});
  localparam [4:0] p13 = (-3'sd2);
  localparam [5:0] p14 = (+((-(3'sd0))!=((-3'sd2)?(3'd5):(5'd6))));
  localparam signed [3:0] p15 = {(-{(+((-5'sd11)?(4'd4):(2'd1))),(-((-5'sd0)&&(4'd8))),(~((-5'sd10)&(5'sd11)))})};
  localparam signed [4:0] p16 = (3'sd3);
  localparam signed [5:0] p17 = (~|(3'sd2));

  assign y0 = ($unsigned(((p3?b1:b2)>$unsigned($signed((b1^~a4))))));
  assign y1 = (b1^p17);
  assign y2 = ((&((p0==p16)&(p5>>b0)))>>((p1^~p3)^~(p5<=p3)));
  assign y3 = {1{((((&p15)<={1{b0}})<<<$unsigned((a4!=a3)))||{4{(p6^~p3)}})}};
  assign y4 = (~&((a3?p15:b4)?((~b4)||(5'd19)):((3'sd1)==(b1%b1))));
  assign y5 = ((a1<<p15)^(b2===a0));
  assign y6 = ($signed(((+b3)<={3{b5}}))&(-5'sd12));
  assign y7 = ({(a2!=p10),(4'd0),{b0,p3}}|(-3'sd1));
  assign y8 = (((p4?p1:p2))?{(p6?p2:b5)}:{{a4},(p7),{p12,p17,p5}});
  assign y9 = {2{(6'd2 * (2'd0))}};
  assign y10 = (+((~^(-a1))<<(b1^b2)));
  assign y11 = {{1{{4{a5}}}},(a3>=b3)};
  assign y12 = (!(~(^(~|(^(~|(~(+(-(|(~p14)))))))))));
  assign y13 = ((+b2));
  assign y14 = ((((b4)?(b3?b0:a5):$unsigned(p6))?$unsigned(($signed(b0)?(a4?p3:b0):(p4))):($signed(p10)?$signed(b1):(b4?p4:p5))));
  assign y15 = (2'd1);
  assign y16 = {4{b3}};
  assign y17 = {(b1>>>p6),(~p14)};
endmodule
