module expression_00323(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(4'sd1)}};
  localparam [4:0] p1 = (((2'sd1)?(5'sd10):(-3'sd2))/(-2'sd0));
  localparam [5:0] p2 = ((3'd0)?(5'sd8):(2'd2));
  localparam signed [3:0] p3 = (((3'd7)+(2'sd0))!=((5'd26)>=(-3'sd1)));
  localparam signed [4:0] p4 = (-3'sd2);
  localparam signed [5:0] p5 = (3'd3);
  localparam [3:0] p6 = (+((-3'sd0)||(2'sd0)));
  localparam [4:0] p7 = (~&(+{2{{3{(-3'sd0)}}}}));
  localparam [5:0] p8 = (-5'sd6);
  localparam signed [3:0] p9 = (-2'sd1);
  localparam signed [4:0] p10 = ((3'd6)^~(2'd3));
  localparam signed [5:0] p11 = ((3'd1)?(5'd31):(4'sd7));
  localparam [3:0] p12 = (+({2{((-5'sd10)<<<(3'd6))}}|(((5'sd3)>=(3'sd2))|(-((5'd25)==(-3'sd0))))));
  localparam [4:0] p13 = (~^(~^(((-2'sd0)?(3'd3):(4'd10))?(&(5'd2)):(-(2'sd0)))));
  localparam [5:0] p14 = (((3'd3)?(2'd2):(4'sd1))>>>{(-2'sd1)});
  localparam signed [3:0] p15 = (~|(-4'sd7));
  localparam signed [4:0] p16 = (&(&(2'sd0)));
  localparam signed [5:0] p17 = (!{(^{4{(-5'sd7)}}),(~(&((^(4'd0))^{(5'd1),(3'sd2)})))});

  assign y0 = ({1{((p8-p10)==(p15<p5))}}<(5'd10));
  assign y1 = (|(((3'sd3)<=(-(p2?p6:b2)))>>>(2'sd0)));
  assign y2 = $unsigned($signed((5'd2 * $unsigned((b1)))));
  assign y3 = (&((2'sd0)<(~^(~|((5'd28)<=(b5^~a0))))));
  assign y4 = (-5'sd11);
  assign y5 = (((p10<<<a2)?{p10,p1}:(p5<=p10))<=({p2,p14,p15}||(p0<=p2)));
  assign y6 = ({3{(b3&a3)}});
  assign y7 = (b3^a1);
  assign y8 = (3'd1);
  assign y9 = (~(~((p6?p13:p17)?(p6||b0):{p5,b1,b1})));
  assign y10 = {1{{2{(+{3{(~|p9)}})}}}};
  assign y11 = {((p12?p5:a3)?(~^p1):(!p13)),((3'd3)>>(a3?b0:b5)),((p11-a0)|(4'd2 * b0))};
  assign y12 = {(+({{b4,b0},{a0,a4}}-{$unsigned({{a0,a2,b3},{4{a2}}})}))};
  assign y13 = ((p12?p8:b5)?(p4?p16:p10):(4'd2));
  assign y14 = (4'd11);
  assign y15 = (($signed(((~^$signed(b4)))))<<((p6?b3:p17)?(a1?p5:p13):(p15)));
  assign y16 = ({3{(a3===b3)}}>>(((p1>>>b0)|{1{a5}})<<<(6'd2 * (3'd6))));
  assign y17 = (4'd2);
endmodule
