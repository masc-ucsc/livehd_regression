module expression_00124(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(~|{1{(!{(-5'sd4),(2'd1),(-5'sd4)})}}));
  localparam [4:0] p1 = ((((4'sd4)<=(5'd6))===((5'd16)>=(2'sd0)))&&(((3'd6)!==(5'd8))>=((-4'sd7)^(2'sd0))));
  localparam [5:0] p2 = {3{((2'd0)?(2'd2):(-2'sd1))}};
  localparam signed [3:0] p3 = ((&(5'd2))&&((4'd9)>>>(-3'sd3)));
  localparam signed [4:0] p4 = (~|(^{2{(4'sd3)}}));
  localparam signed [5:0] p5 = ((|((5'sd7)>>>(4'sd7)))>>>(((4'd11)?(5'd26):(-4'sd5))>>>((5'd28)?(5'd5):(4'd14))));
  localparam [3:0] p6 = ((|((-2'sd0)&(-5'sd9)))?(3'd1):(4'd2 * ((4'd5)?(3'd1):(3'd7))));
  localparam [4:0] p7 = (3'sd3);
  localparam [5:0] p8 = {(!((~|(((3'd2)+(2'd0))+(~&(2'sd0))))>={((2'd1)&(4'sd5)),((5'sd6)||(4'd0))}))};
  localparam signed [3:0] p9 = ((3'd7)?(5'd16):(-2'sd0));
  localparam signed [4:0] p10 = (-((~(|(-4'sd1)))/(-4'sd6)));
  localparam signed [5:0] p11 = ((!(((5'd9)+(2'd0))<((4'd11)*(3'd5))))===(^(!(~&(&(^((5'sd7)^(-4'sd7))))))));
  localparam [3:0] p12 = (~&(2'd2));
  localparam [4:0] p13 = {({((-3'sd3)?(4'd8):(4'd10))}?{(5'd10),(-4'sd1),(5'sd0)}:{(5'd8),(5'd8),(3'sd2)})};
  localparam [5:0] p14 = {3{(5'sd5)}};
  localparam signed [3:0] p15 = {2{(-3'sd2)}};
  localparam signed [4:0] p16 = {(3'sd2),(5'd1),(2'd3)};
  localparam signed [5:0] p17 = ({4{(-5'sd11)}}<=(4'd2 * (3'd5)));

  assign y0 = {3{p8}};
  assign y1 = {((-4'sd4)&{4{a1}})};
  assign y2 = (b5!==b2);
  assign y3 = ({3{{p10,b1}}}^~($signed((p9<a1))?{1{(a2-p15)}}:(a2?p16:a2)));
  assign y4 = $unsigned({p14,p15,p0});
  assign y5 = {1{(3'd2)}};
  assign y6 = ((~^(~($signed(b4)<<<(p8||p4))))<<<$unsigned(((p6)>>$unsigned(p4))));
  assign y7 = (2'd3);
  assign y8 = ((+(5'd17))&{b0,b3,a2});
  assign y9 = {4{b2}};
  assign y10 = (2'd3);
  assign y11 = ({3{a0}}?((a1?a0:b4)===(a5?a5:b2)):(b2?a1:p12));
  assign y12 = ({a0}==$unsigned(a4));
  assign y13 = (p13<<<p17);
  assign y14 = ((p16?p14:a1)?$signed(p16):(p7?p4:p12));
  assign y15 = (3'd0);
  assign y16 = (4'd4);
  assign y17 = (((+(4'd2))>=(-(-4'sd3)))?(~((a2!=b0)?(a0>>b2):(b1?p5:a2))):((p16<a3)<<(^{2{b1}})));
endmodule
