module expression_00197(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{1{(4'd12)}},(-2'sd1)};
  localparam [4:0] p1 = (~((-2'sd0)?(-2'sd0):(-3'sd1)));
  localparam [5:0] p2 = (5'd21);
  localparam signed [3:0] p3 = (({{(2'sd0),(5'd0),(2'sd0)}}=={(-3'sd3),(2'd0),(-5'sd2)})<=(+(-3'sd1)));
  localparam signed [4:0] p4 = (!(~&(-{2{{2{{3{(3'sd2)}}}}}})));
  localparam signed [5:0] p5 = (((~&(+(-4'sd3)))>>((2'd0)?(3'd7):(2'sd0)))^~(((2'd2)<(5'd29))>>(^((2'sd1)>>(3'd6)))));
  localparam [3:0] p6 = ((({4{(3'd6)}}!==((-5'sd14)>=(4'd13)))^~(4'sd6))!==(5'sd14));
  localparam [4:0] p7 = (+(|((3'd4)?(3'd7):(2'd3))));
  localparam [5:0] p8 = (3'd1);
  localparam signed [3:0] p9 = ((3'sd3)==(-4'sd7));
  localparam signed [4:0] p10 = (&({{(4'd3),(3'd0),(5'sd14)}}<=((-5'sd0)<<(3'sd2))));
  localparam signed [5:0] p11 = ((4'sd3)^~(2'd3));
  localparam [3:0] p12 = {3{((2'sd1)?(-3'sd0):(5'd2))}};
  localparam [4:0] p13 = (-2'sd0);
  localparam [5:0] p14 = {{(2'sd1),(5'd13),(3'd7)},({4{(2'd0)}}!={1{(5'd24)}}),({3{(2'd2)}}!==((5'sd3)||(5'sd8)))};
  localparam signed [3:0] p15 = (-(((5'd2)?(4'd10):(3'sd2))?(~&((-3'sd2)?(2'd2):(3'd3))):(~&((-3'sd0)^~(4'd3)))));
  localparam signed [4:0] p16 = ((4'sd3)>>(((5'd10)>=(2'd2))?(5'd3):(-3'sd3)));
  localparam signed [5:0] p17 = {(~(-4'sd7)),((-4'sd2)!=(2'd2)),{(-5'sd2),(4'd10),(5'd22)}};

  assign y0 = ((p2<=p1)<(6'd2 * p7));
  assign y1 = (~&((~&a2)?(a0%a1):(-a1)));
  assign y2 = (2'sd0);
  assign y3 = ((|((p6&&p14)>>(p15?p1:p16)))?{{2{{4{p9}}}}}:({b4,a5}==={a0,a4}));
  assign y4 = ((~((b1==p7)<<(p4?p0:a3)))?(5'sd3):(~^(&((-3'sd2)?(b1^~p10):(~^p2)))));
  assign y5 = (2'sd0);
  assign y6 = (~|((p11?p5:b4)?(~(~(~|p5))):(b0?a5:a5)));
  assign y7 = $unsigned((~^{(+(2'd2)),(^(+(|(~^b3))))}));
  assign y8 = ({3{(b4&&a2)}}^({1{{4{b5}}}}==((a5==a3)<{2{b4}})));
  assign y9 = $signed((p1>=p9));
  assign y10 = ((~((6'd2 * p2)%a2))>=((~^((~a3)<(p8-b3)))<<(~|((p2^b2)&&(p7<<p2)))));
  assign y11 = (p3?a0:p1);
  assign y12 = (&{3{(&(!p4))}});
  assign y13 = (^{4{(a5^~b3)}});
  assign y14 = {3{$unsigned((+{2{a0}}))}};
  assign y15 = {4{(b2!==a4)}};
  assign y16 = {2{{(-(~(2'sd1)))}}};
  assign y17 = ((b1<<<b4)?(a2?a3:a2):(b5===a1));
endmodule
