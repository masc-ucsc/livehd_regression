module expression_00332(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(-2'sd0),(3'd6),(2'd0)}^~((5'sd12)?(4'sd5):(4'd10)));
  localparam [4:0] p1 = ((3'd4)&&(3'd2));
  localparam [5:0] p2 = ((((-3'sd3)?(3'd0):(-2'sd0))-((-2'sd1)>(-3'sd2)))?(((3'd1)&(5'sd13))>>>((2'sd0)?(5'd13):(4'sd1))):((2'd1)?(2'd1):(2'sd0)));
  localparam signed [3:0] p3 = (~{4{(~|((5'sd5)<<(3'sd2)))}});
  localparam signed [4:0] p4 = {3{(-3'sd1)}};
  localparam signed [5:0] p5 = (-5'sd14);
  localparam [3:0] p6 = (|(5'd2 * (2'd2)));
  localparam [4:0] p7 = ((~&(3'd1))<<(3'd7));
  localparam [5:0] p8 = {{4{{4{(5'd27)}}}}};
  localparam signed [3:0] p9 = {4{((2'd3)===(2'sd0))}};
  localparam signed [4:0] p10 = (((^(5'd15))||{3{(2'd3)}})?((4'd2)?(-5'sd5):(-5'sd2)):(((2'd0)+(2'sd0))>>{4{(2'sd0)}}));
  localparam signed [5:0] p11 = (((-4'sd0)?(5'd25):(5'd28))?((2'sd0)?(3'd2):(5'd5)):((2'd1)<<<(3'sd0)));
  localparam [3:0] p12 = (!(5'sd8));
  localparam [4:0] p13 = ((~{(-3'sd2)})?(2'd1):{4{(-3'sd3)}});
  localparam [5:0] p14 = (^((((5'd30)-(2'sd0))||((-5'sd0)<(-5'sd10)))!={(~|(5'd2 * ((2'd1)&(4'd15))))}));
  localparam signed [3:0] p15 = {((~^(2'd0))||{(~^(2'sd1))}),({(2'd3),(2'd3)}^{(2'd1),(4'd4),(4'd3)})};
  localparam signed [4:0] p16 = ({((5'd31)<<(5'd7)),(4'd2 * (2'd0))}>>>(((-5'sd0)+(-4'sd4))^~((5'd8)>(3'd5))));
  localparam signed [5:0] p17 = (+(^(^(~|((~^(-(4'd12)))?((5'sd0)^(5'sd3)):(~|(|(-2'sd1))))))));

  assign y0 = (~|(p0?p5:p1));
  assign y1 = {{2{b2}}};
  assign y2 = ((|((p3<=a0)>=(|(!p12))))==((!(!(2'd0)))<(&(a0<=p14))));
  assign y3 = (-5'sd13);
  assign y4 = ((((b3)?(&a4):{a0,p10}))<($signed((+b2))?(a4===b0):{$signed(p5)}));
  assign y5 = ((p11)>>>$signed(p4));
  assign y6 = (!a4);
  assign y7 = ((p2?p3:p12)?(p12?p7:a2):(p15?p0:p16));
  assign y8 = (~&(-2'sd1));
  assign y9 = ((a5+p7)/p5);
  assign y10 = (~(~^b5));
  assign y11 = {(((3'sd1)?(p4?p6:p13):(6'd2 * p8))&({(2'd3)}<<{p3,p12,p8}))};
  assign y12 = ((p15>>p4)>=(p3>p12));
  assign y13 = (!(~|(~^((p4&b0)>=(~p6)))));
  assign y14 = (-4'sd2);
  assign y15 = (^((|((^(~&(!a2)))^~((a4^a5)<<(b3>=b4))))|(-4'sd1)));
  assign y16 = ($unsigned((!b0))%a2);
  assign y17 = (((4'd9)|((5'd2 * p2)||(b4?b3:a0)))||((4'd3)?(4'd0):{a2,a1,a2}));
endmodule
