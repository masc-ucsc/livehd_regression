module expression_00285(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(6'd2 * ((4'd6)>=(2'd2))));
  localparam [4:0] p1 = ({(-2'sd0),{(-3'sd0),(-2'sd0)}}^~(^(^(4'd13))));
  localparam [5:0] p2 = (+((((4'd15)<(-2'sd0))-((5'sd5)!=(-4'sd3)))?(&((-2'sd0)&&(-2'sd0))):(!((-5'sd1)>>>(3'd0)))));
  localparam signed [3:0] p3 = (({4{(5'sd7)}}?((4'sd2)>(4'd2)):((4'd4)?(2'd0):(2'sd0)))&(|(((-2'sd0)|(3'd0))!=(&(4'sd7)))));
  localparam signed [4:0] p4 = (-4'sd7);
  localparam signed [5:0] p5 = ((-5'sd0)?(5'sd7):(5'sd15));
  localparam [3:0] p6 = ((((2'd0)>>(5'd6))+((5'sd3)^(4'd12)))>(4'd2 * (5'd2 * (2'd3))));
  localparam [4:0] p7 = (3'd6);
  localparam [5:0] p8 = (&(~|((&(3'd2))>((2'sd0)>=(-4'sd1)))));
  localparam signed [3:0] p9 = (((4'sd6)<=(-5'sd1))?(~&((-2'sd0)*(-5'sd1))):((2'sd1)?(-2'sd0):(3'd1)));
  localparam signed [4:0] p10 = (4'd2 * (2'd1));
  localparam signed [5:0] p11 = ({1{{4{(-3'sd2)}}}}+{3{(5'sd12)}});
  localparam [3:0] p12 = (&{2{(5'sd4)}});
  localparam [4:0] p13 = ({1{((-2'sd1)?(-2'sd0):(2'd3))}}?(~^(-4'sd0)):(-5'sd0));
  localparam [5:0] p14 = {2{(5'd25)}};
  localparam signed [3:0] p15 = (~^(^(((-{3{(4'd14)}})!==((5'd26)&(5'd18)))<<(-(~(~^((5'd1)<<<(5'd3))))))));
  localparam signed [4:0] p16 = ((5'sd1)+((((5'd7)>=(-3'sd0))===((2'd1)^~(-3'sd1)))&&({4{(-3'sd2)}}<<(2'sd1))));
  localparam signed [5:0] p17 = (^(+(&(((-4'sd2)?(4'sd2):(5'sd2))^~((3'sd1)<=(-5'sd14))))));

  assign y0 = (~({(b2>a2),(3'sd2),{b5,p0}}>>>{(+b0),{b0,a4},{p7,a2,b4}}));
  assign y1 = {((2'd3)>={b2,a3,p6}),((+p3)-(p13^p9)),(5'd15)};
  assign y2 = (~^((~&(((~|(^(-(|$signed(p5))))))&&(~^(+(~^((|a3)>=(~b5)))))))));
  assign y3 = (^(|{3{{4{p2}}}}));
  assign y4 = ($unsigned($signed((^((2'd3)?(p15>=p9):(p7>=a3))))));
  assign y5 = {{{p12,p0,p17},{(!{p3,p7,p12})}}};
  assign y6 = ((b1?a1:a2)?(b4?a5:b3):(b2?a2:p13));
  assign y7 = (-4'sd6);
  assign y8 = ((4'd11)>(5'sd2));
  assign y9 = (({b5,b4,b0}?(b4?a3:b1):((b3>>>a0)))|{(b0?b0:a4),(a0+a3),$unsigned({b1,a0})});
  assign y10 = (~&(!(-a1)));
  assign y11 = (4'd2 * {a0,p2,p0});
  assign y12 = (p10?p15:p6);
  assign y13 = {(^(~&p1)),(a5!=p12)};
  assign y14 = (~^(5'd2 * (a1>b0)));
  assign y15 = (^{(~(+$unsigned(b2))),(+(|(~b1))),(p11?p11:b4)});
  assign y16 = ((5'd2 * a1)!==(~^(5'd2 * a2)));
  assign y17 = {(a5?p10:p3),(a5?a1:p13),{p7,b3,p5}};
endmodule
