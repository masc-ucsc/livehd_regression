module expression_00167(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd4)/(5'd25))<<<((4'd9)^~(4'd8)))>>((~|(~|(3'd7)))>((2'd2)&(4'd14))));
  localparam [4:0] p1 = (~|(({2{(-4'sd1)}}<<<((3'd0)==(-5'sd11)))<<{(~(5'd16)),(~&(2'd0)),((-2'sd0)&(3'sd0))}));
  localparam [5:0] p2 = ({((3'sd0)>(-5'sd15)),((5'd24)^(-5'sd8)),((-2'sd0)-(2'd3))}>>>{{{(3'sd0),(5'sd10),(4'd0)}},((2'd3)^~(2'd3))});
  localparam signed [3:0] p3 = ({3{(4'sd2)}}?((5'd2 * (2'd1))-((-2'sd1)?(5'd18):(5'd2))):(-((4'd0)<<<(5'd6))));
  localparam signed [4:0] p4 = {(!(-((3'd6)==(5'sd5)))),{{(3'd4)},((-2'sd0)>=(5'd22)),((-4'sd5)<(-4'sd4))}};
  localparam signed [5:0] p5 = {2{(~({1{(3'sd1)}}&&(~&(2'd0))))}};
  localparam [3:0] p6 = (5'd4);
  localparam [4:0] p7 = {4{((4'd9)<(-2'sd1))}};
  localparam [5:0] p8 = (((4'd6)?(2'sd1):(4'sd4))!=={2{(3'd3)}});
  localparam signed [3:0] p9 = {{4{{{1{(4'd10)}}}}}};
  localparam signed [4:0] p10 = {(((3'd3)?(2'sd0):(4'd7))?((3'sd3)>=(4'd2)):{(4'd4)}),(((4'd15)===(-5'sd12))===((3'sd3)&(3'sd1))),{4{(2'd3)}}};
  localparam signed [5:0] p11 = (6'd2 * (~&(5'd23)));
  localparam [3:0] p12 = ((((4'd4)?(-4'sd1):(-4'sd3))&{(3'd5),(2'sd0)})<<(((2'd1)||(2'sd1))^{(-(3'd4))}));
  localparam [4:0] p13 = ((3'd0)^(2'd0));
  localparam [5:0] p14 = (2'd2);
  localparam signed [3:0] p15 = ({4{(2'sd1)}}?((2'd2)?(4'sd3):(5'd4)):(2'd0));
  localparam signed [4:0] p16 = {{(5'd31),(3'd6),(-3'sd0)},{(5'sd13),(-2'sd1)},{(3'sd2),(4'd13),(4'd12)}};
  localparam signed [5:0] p17 = {({(2'd3),(5'sd14),(2'd0)}!==((2'sd0)<<(-4'sd1))),(^({(5'd23),(3'd7),(3'd0)}>>>(~&(2'd1)))),(((2'd3)-(-4'sd1))==(^(5'd27)))};

  assign y0 = {({p5,p13,p13}?(-(p11?p3:p7)):(4'sd2)),(4'sd7)};
  assign y1 = {(p4<=b4),(p17>>p10)};
  assign y2 = {1{(~|{{2{a1}},{1{{b0,a2,p6}}}})}};
  assign y3 = $unsigned({{(~p14),{a4,b3}},(+({b0,p15,p0}+(b1==p1))),((+$unsigned($unsigned(a2))))});
  assign y4 = ((3'd7)<<<(~|(4'sd7)));
  assign y5 = (((~p0)?(p7?p2:p15):(b3?p9:b5))?(!(~&(+(a5?p3:b5)))):{(b1>b0),(~&a1),(~&b5)});
  assign y6 = (!(&(((~|p2)%p16)^(~^(~^(p10))))));
  assign y7 = (((a1?p15:b5)?(~^p17):(p4?p13:p0))?(!(~(|(p0?p2:p16)))):(~|((p12?a1:p17)?(p3?p13:p6):(a4?b5:a5))));
  assign y8 = (~^(~|p12));
  assign y9 = (&(((a0?b0:a3)<<(&(a0||a4)))||(((p7?a0:b3)?(a2?b1:a2):$unsigned(a1)))));
  assign y10 = {3{{3{{1{p15}}}}}};
  assign y11 = (a5?a4:a3);
  assign y12 = (5'd10);
  assign y13 = ((3'd1)>={((2'd1)&((b4&&a3)>>{4{b5}}))});
  assign y14 = {p1,p4,b4};
  assign y15 = (p4?p17:p11);
  assign y16 = (~|(!((!(4'd2 * p0))?(&(b1+b2)):((-4'sd6)>>$unsigned(a5)))));
  assign y17 = ((|(~^((a1!=b2)&&{3{p8}})))&&(^((p1+p13)<=(p0<<<b2))));
endmodule
