module expression_00867(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(4'd4));
  localparam [4:0] p1 = ({{(5'd20),(2'd0)},{4{(-3'sd1)}}}>>(~^(^(~^(-4'sd6)))));
  localparam [5:0] p2 = (-{2{(-((5'd3)|(2'sd1)))}});
  localparam signed [3:0] p3 = (2'd2);
  localparam signed [4:0] p4 = (5'd20);
  localparam signed [5:0] p5 = (~|((~((3'sd1)?(4'd15):(2'sd0)))?(!{{1{(2'd3)}}}):({1{(3'd0)}}^(|(-5'sd7)))));
  localparam [3:0] p6 = ((^(((2'd1)>=(-2'sd1))?{3{(5'd11)}}:((5'd14)!==(2'sd0))))^({1{{4{(-2'sd0)}}}}|{1{((5'd5)<<<(5'd29))}}));
  localparam [4:0] p7 = ({1{((2'sd0)?(5'sd8):(-4'sd4))}}?(5'd2 * {(3'd5),(5'd4)}):{(~(6'd2 * (4'd4)))});
  localparam [5:0] p8 = (~^((3'd7)?(5'sd12):(2'd3)));
  localparam signed [3:0] p9 = (((2'd3)>=(-5'sd1))&&(&(5'd2 * (3'd0))));
  localparam signed [4:0] p10 = (-4'sd5);
  localparam signed [5:0] p11 = {3{{4{(3'd4)}}}};
  localparam [3:0] p12 = {1{{1{(3'sd1)}}}};
  localparam [4:0] p13 = (5'd2 * ((4'd10)==(2'd2)));
  localparam [5:0] p14 = (-(((4'sd1)||(-4'sd2))*(~^(4'd9))));
  localparam signed [3:0] p15 = (^{1{(5'd25)}});
  localparam signed [4:0] p16 = {{{2{(4'd14)}},{(2'sd0)},{(5'sd2),(4'd7),(4'd0)}},{{(4'd2),(5'd15)},{(5'd29)},{3{(-3'sd2)}}}};
  localparam signed [5:0] p17 = (3'sd1);

  assign y0 = (~((~&(~(&b0)))&&(~&(b5===b3))));
  assign y1 = {1{b2}};
  assign y2 = {1{{3{(a5^~p14)}}}};
  assign y3 = ({{($signed((~&b1)))}}!==(-$unsigned({a1,a0,b2})));
  assign y4 = (5'sd6);
  assign y5 = (({1{p0}}>>{a5,p14}));
  assign y6 = {(((p4)?{a0,a0}:{4{p9}})?{4{a3}}:((|a4)?(a3>=b2):(p8)))};
  assign y7 = ($signed($signed((~$unsigned(((b5<<<b3)<(^p10))))))-((b1?a5:b1)===(b2?a1:a2)));
  assign y8 = {4{b2}};
  assign y9 = $signed((~^(!(~&(!$unsigned({3{(&(p16?p15:p10))}}))))));
  assign y10 = ((5'd3)<=(^(-4'sd5)));
  assign y11 = {2{(((p5?p3:p0)==(p15+p15))!=((p2?p8:p14)?{1{p0}}:(2'd0)))}};
  assign y12 = (((a2==p6)/b5)-(((a2^a5))===(b0>>b1)));
  assign y13 = $signed((-5'sd9));
  assign y14 = ((p9>>>p15)!=(p15<=b0));
  assign y15 = (((p0||a0)^(-5'sd2))^(4'd13));
  assign y16 = ((a0?p13:b0)>>{3{a4}});
  assign y17 = (b4!=b4);
endmodule
