module expression_00179(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(-2'sd0)}>{(3'd7),(2'd3)});
  localparam [4:0] p1 = (4'sd4);
  localparam [5:0] p2 = {3{((2'sd0)||((3'sd0)<(4'd8)))}};
  localparam signed [3:0] p3 = {2{((5'd29)?((-2'sd1)!==(3'd7)):((4'd3)<=(2'd1)))}};
  localparam signed [4:0] p4 = (+(~^((~&(~&((4'sd4)?(4'sd3):(4'd6))))?(((3'sd2)?(5'd23):(-5'sd15))&&((5'sd8)?(2'd3):(4'sd2))):((3'sd3)?(5'sd10):(2'sd1)))));
  localparam signed [5:0] p5 = ((-4'sd6)?(~|(&((3'd3)?(5'sd0):(3'd1)))):(-(((-4'sd7)>(2'd1))^~{2{(-5'sd5)}})));
  localparam [3:0] p6 = {2{(((-5'sd12)>(3'd6))&&(~|(-4'sd1)))}};
  localparam [4:0] p7 = ((!(~|((-3'sd2)!=(2'd0))))>>((~|(3'd4))<=((4'sd3)>(2'sd1))));
  localparam [5:0] p8 = (-(&(-2'sd0)));
  localparam signed [3:0] p9 = (5'd16);
  localparam signed [4:0] p10 = ((5'd21)?(4'sd5):(4'd0));
  localparam signed [5:0] p11 = (&(-2'sd0));
  localparam [3:0] p12 = (!(+(4'd2 * (5'd29))));
  localparam [4:0] p13 = (3'd2);
  localparam [5:0] p14 = (!((3'sd0)<<(4'd5)));
  localparam signed [3:0] p15 = (((3'sd0)^(4'd11))?(-{4{(5'd0)}}):(5'd2 * (5'd0)));
  localparam signed [4:0] p16 = (^(5'sd9));
  localparam signed [5:0] p17 = ((((3'd2)===(3'd2))>>((5'sd9)/(3'd1)))?(((3'sd2)?(2'd3):(3'd0))?((-3'sd1)!=(2'sd0)):((-4'sd0)^~(2'd1))):(((5'd9)?(3'd6):(4'sd0))&&((2'sd1)?(-3'sd1):(4'sd0))));

  assign y0 = {(a0?a5:p17),(2'd3),{1{{3{a2}}}}};
  assign y1 = {4{b0}};
  assign y2 = {1{{4{(^{2{{a2,b4,a0}}})}}}};
  assign y3 = {{(p3+b0),{b1,b3,b4}}};
  assign y4 = {2{((~^(!p16))+{1{{4{p8}}}})}};
  assign y5 = (|p11);
  assign y6 = {2{$signed({b1,b0})}};
  assign y7 = (-(~&(~^(&($unsigned($signed((p15/b3))))))));
  assign y8 = ((p1?b3:a2)^~(a1?a0:p3));
  assign y9 = (a0|p0);
  assign y10 = (~|{((|(b1===a2))<={(~&p12)}),((p7==a3)?(5'd3):(a0?a3:p2)),(4'd11)});
  assign y11 = {1{(!{{4{p7}},(|a4)})}};
  assign y12 = (({b0,p8,a2}?(&p12):(~|p10))?{(|(~(a1?b0:a3)))}:({2{p9}}?(p4?p0:p7):{1{p5}}));
  assign y13 = (((~&p4)+(-4'sd7))<=$unsigned((+(p10-p10))));
  assign y14 = ($signed(p1)!=(p12||p5));
  assign y15 = (|({{4{b2}}}>>>{1{{(&(a2?b2:p0))}}}));
  assign y16 = ((|(^b0))%b3);
  assign y17 = (((b0)?{b2,b0}:{b2,b5})?((a5)?(&a3):(a3^b3)):($unsigned({a4})&{a2,a4,a3}));
endmodule
