module expression_00367(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'd28)||(~^(4'd4)))<(~(~|((-2'sd0)>>>(-5'sd2)))));
  localparam [4:0] p1 = (!(((~|(4'd6))?((-4'sd1)?(2'd0):(-5'sd8)):((5'sd2)?(-3'sd1):(5'd18)))!==(~(~^((2'sd1)?(-5'sd2):(4'd5))))));
  localparam [5:0] p2 = (|{(4'd13),(5'd13)});
  localparam signed [3:0] p3 = ((4'd1)<<(3'd0));
  localparam signed [4:0] p4 = ((~((&(4'd4))<=((-3'sd2)?(3'd1):(4'd2))))?(&((^(-3'sd3))>=((-2'sd1)?(-2'sd0):(-2'sd1)))):(~&(^(&(~^(4'd15))))));
  localparam signed [5:0] p5 = (-((((-5'sd10)?(5'sd3):(-5'sd9))?{4{(-5'sd4)}}:{4{(2'd2)}})^(+(~^(~((4'd11)?(-4'sd2):(3'd7)))))));
  localparam [3:0] p6 = (((4'd13)>>>(-5'sd11))===((-4'sd4)<=(5'd7)));
  localparam [4:0] p7 = ((2'sd1)^(2'sd0));
  localparam [5:0] p8 = ((((2'd1)<<(3'sd3))<((3'd5)===(2'sd0)))>>>(~|(~(3'd6))));
  localparam signed [3:0] p9 = (-5'sd0);
  localparam signed [4:0] p10 = (!({1{(4'd6)}}?((4'd2)<(2'd1)):(5'd2 * (5'd26))));
  localparam signed [5:0] p11 = {4{(2'd0)}};
  localparam [3:0] p12 = ((-(~^(4'd3)))<<(6'd2 * (4'd10)));
  localparam [4:0] p13 = {(((4'sd0)<(2'd3))>>>((3'd6)!==(5'd29))),(((5'd6)===(2'sd0))^~{2{(5'd16)}})};
  localparam [5:0] p14 = (~|(((-5'sd15)>(2'd2))!=((4'sd5)<<<(3'd6))));
  localparam signed [3:0] p15 = ({{(5'd19),(-4'sd6)},{3{(4'sd0)}},{1{(2'd3)}}}>>{4{{(5'd13)}}});
  localparam signed [4:0] p16 = ((+(4'sd6))?((2'd1)^~(2'd0)):(!(3'd5)));
  localparam signed [5:0] p17 = ((((4'sd5)-(-3'sd1))&&((-4'sd3)<=(-3'sd2)))<<(((4'd13)>=(-2'sd0))%(3'd4)));

  assign y0 = ((a4?a3:b2)-(p9<<a3));
  assign y1 = (3'd0);
  assign y2 = ($signed((a1===a2)));
  assign y3 = (-((^(a3<<b0))||({1{p5}}<<<(~^p1))));
  assign y4 = ((p11^a3)>=$signed((b4)));
  assign y5 = {3{{4{p16}}}};
  assign y6 = (((b1?a5:b1)^~(b5|b4))===((a4?b3:a5)|(a0^a3)));
  assign y7 = (~^(&(4'sd3)));
  assign y8 = ((~|((5'd2 * p13)^{p13,b4,a2}))+((-b5)-(|a0)));
  assign y9 = (|(5'd21));
  assign y10 = ((!(-4'sd7))>>>{3{p0}});
  assign y11 = $signed(b5);
  assign y12 = $signed((!(5'd20)));
  assign y13 = ({{b3,b4,p4}}>((b2|b2)>(b4?a0:b3)));
  assign y14 = ({$signed({($unsigned(p15)),{a0,p12,p12}})}|$unsigned(((4'd14)|{3{a5}})));
  assign y15 = ((b4^~a1)?(b0?p13:p3):(!(b3!=b2)));
  assign y16 = {(~&(|$signed((^p13)))),({(!(p17?p11:p10))}),((p9?p10:p9)?$unsigned(p17):(p0?p2:p8))};
  assign y17 = (~^b4);
endmodule
