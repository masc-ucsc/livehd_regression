module expression_00764(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(((2'd0)==(3'sd3))<<<{(4'sd0),(2'd3),(-4'sd0)})}};
  localparam [4:0] p1 = (5'sd4);
  localparam [5:0] p2 = (({4{(2'sd1)}}?(-3'sd3):((-5'sd0)<=(2'sd1)))<(((4'd12)?(4'sd0):(4'sd5))||((-2'sd0)^~(5'd21))));
  localparam signed [3:0] p3 = (+{{(4'd4),(2'd3),(-2'sd0)}});
  localparam signed [4:0] p4 = (-2'sd1);
  localparam signed [5:0] p5 = {4{{4{(3'sd2)}}}};
  localparam [3:0] p6 = (((3'd7)?(3'd7):(5'd2))?((3'd1)<(3'd1)):((4'sd1)!=(-3'sd2)));
  localparam [4:0] p7 = (~&({1{((5'd4)?(-3'sd3):(4'd9))}}?({3{(5'sd4)}}===(^(2'sd1))):{4{(4'd2)}}));
  localparam [5:0] p8 = (-5'sd11);
  localparam signed [3:0] p9 = ((3'd5)?(2'sd0):(4'd1));
  localparam signed [4:0] p10 = (4'd5);
  localparam signed [5:0] p11 = ((4'd0)<<<(-4'sd1));
  localparam [3:0] p12 = ((^{{(-2'sd1)},((-2'sd1)-(2'd2)),{(2'd2),(3'sd2)}})!==((-((5'd15)===(5'sd14)))>>(|(-(5'sd10)))));
  localparam [4:0] p13 = ((((3'd4)*(5'sd5))?((-4'sd1)>(2'sd1)):((2'd3)?(5'sd10):(4'sd1)))==((6'd2 * (5'd16))?((3'sd3)===(-5'sd0)):((3'd3)?(-4'sd4):(4'd11))));
  localparam [5:0] p14 = {(4'd9)};
  localparam signed [3:0] p15 = (^(~|(4'd12)));
  localparam signed [4:0] p16 = (((5'd24)?(-3'sd2):(5'd26))>>((-5'sd13)/(3'd7)));
  localparam signed [5:0] p17 = {({((2'd3)?(3'd3):(-4'sd6))}?(((-2'sd0)&&(4'd15))^((2'd0)<<<(2'd1))):(5'd2 * ((4'd1)<<<(5'd6))))};

  assign y0 = $unsigned(((p15>=p10)%p10));
  assign y1 = ((!{p12,p4,p15})+((4'd11)^$unsigned(b0)));
  assign y2 = {1{{4{(~|(4'd10))}}}};
  assign y3 = (~^p12);
  assign y4 = (((5'd12)>>>((a2!==b2)<<<(a2*p4)))+((b2>>>p0)%a3));
  assign y5 = {1{({1{(b1&a5)}}^(b3!=b2))}};
  assign y6 = (!$signed(p3));
  assign y7 = $unsigned((p6?b4:b4));
  assign y8 = {a5,p14};
  assign y9 = (p16&p14);
  assign y10 = {4{$signed({4{b2}})}};
  assign y11 = {3{(a0?b0:a1)}};
  assign y12 = (!(~&$signed({3{({3{p14}})}})));
  assign y13 = $signed((3'd4));
  assign y14 = (((!(p7^~b1))|{4{p14}})<<<((&$signed((|((~p8)>>>(-a2)))))));
  assign y15 = (^((p8)||(-4'sd7)));
  assign y16 = (5'd20);
  assign y17 = (b5+b5);
endmodule
