module expression_00665(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((&(&((-3'sd0)<<<(5'd11))))^(~^(~(~(3'd6)))))>>>(((5'd8)?(-5'sd10):(4'd14))^((4'sd5)?(2'sd0):(5'd11))));
  localparam [4:0] p1 = (+(4'sd6));
  localparam [5:0] p2 = ((|((~|(3'sd3))?{(4'sd4),(5'sd10)}:((2'd3)?(3'd6):(4'sd1))))>>>((-((3'sd1)?(4'd6):(2'd3)))>>{{1{(3'd7)}}}));
  localparam signed [3:0] p3 = (4'd14);
  localparam signed [4:0] p4 = ((((3'd7)===(3'd3))?((3'd7)>>>(3'sd2)):(~|(-4'sd0)))<=(((3'd1)<<<(2'sd1))<<<((5'd1)*(3'sd2))));
  localparam signed [5:0] p5 = {(5'd18),(2'sd0)};
  localparam [3:0] p6 = (4'd2 * ((3'd2)*(5'd28)));
  localparam [4:0] p7 = (+(^({(+((-2'sd0)|(5'd12)))}<=(((-4'sd7)!=(2'sd0))-{(3'd1)}))));
  localparam [5:0] p8 = (|(2'd3));
  localparam signed [3:0] p9 = (((3'd6)?(4'sd3):(2'sd0))?(2'd1):((4'd12)?(5'sd15):(5'd14)));
  localparam signed [4:0] p10 = ((~|(2'd2))?((5'd27)===(3'd6)):(|(~|(5'd4))));
  localparam signed [5:0] p11 = ((-3'sd3)>=(4'd9));
  localparam [3:0] p12 = ((~&(^((-(2'sd1))>((3'd3)!==(2'sd0)))))<<(((4'sd2)!=(3'd6))<=((4'd1)>>(3'sd3))));
  localparam [4:0] p13 = (!((^(~(~^(4'd15))))>>({2{(4'sd3)}}<<{2{(5'd7)}})));
  localparam [5:0] p14 = ((4'd3)>>((5'sd8)|((3'd1)>>(3'd1))));
  localparam signed [3:0] p15 = (3'd4);
  localparam signed [4:0] p16 = (3'd2);
  localparam signed [5:0] p17 = (((4'sd0)&&(-5'sd10))/(2'sd0));

  assign y0 = {{((b1)||(p14>a3))},(!$signed($unsigned((~^(3'd3)))))};
  assign y1 = (+{(~&({{b2}}>>{b3,b2})),{({p16}?(p3>=a5):(a3<<<b2))}});
  assign y2 = (($signed((3'd3))<<($signed(a3)|(b0&&a1)))!==((-4'sd4)));
  assign y3 = {(a3&p9),{(a1&b5)}};
  assign y4 = (b3&&p2);
  assign y5 = {$unsigned($unsigned((&{1{({1{({p12,p11,p3})}})}})))};
  assign y6 = ({2{{3{b0}}}}?((a4>b3)>>>{4{b5}}):{2{(&(a5?a2:a5))}});
  assign y7 = (~((^({4{a0}}<<(b3?b1:p11)))?(~&(p1?a4:p3)):{(b0?p7:p5),(a0?a3:p5)}));
  assign y8 = ((p0==p17)>>{4{a2}});
  assign y9 = (!p15);
  assign y10 = {2{{4{(|b0)}}}};
  assign y11 = (5'sd13);
  assign y12 = (+(-4'sd1));
  assign y13 = ({3{(a1||b1)}}?((p12?b5:p10)?(&a3):(a1^a0)):({4{p9}}>>(b2!==a2)));
  assign y14 = ((b5&&a3)!=(b1!==b4));
  assign y15 = (((~(a4>p8))<<((b3+a4)|(4'd5)))<=(3'd6));
  assign y16 = ((&$signed($unsigned((!(-$signed(($unsigned({1{({2{{3{(+p10)}}}})}})))))))));
  assign y17 = (4'd5);
endmodule
