module expression_00992(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{((4'sd3)||(-5'sd14))}};
  localparam [4:0] p1 = ((2'd1)+(+{4{(-4'sd0)}}));
  localparam [5:0] p2 = (-2'sd0);
  localparam signed [3:0] p3 = {(-5'sd14),{2{(5'sd5)}},(((4'd9)>=(3'd2))?((5'd23)+(-3'sd3)):(-2'sd1))};
  localparam signed [4:0] p4 = ((((5'd12)>=(-4'sd4))==(!(-4'sd7)))&({(2'sd0)}<<((5'sd14)!==(5'd23))));
  localparam signed [5:0] p5 = (2'sd1);
  localparam [3:0] p6 = {2{((4'sd2)?(-4'sd0):(4'd3))}};
  localparam [4:0] p7 = (~^(-(((2'd1)?(2'sd0):(3'sd1))?((4'sd6)?(4'sd2):(-5'sd5)):{(2'd3),(2'sd1),(-2'sd1)})));
  localparam [5:0] p8 = {1{(+(((5'sd14)?(3'sd1):(3'sd3))>>(~&((5'sd10)==(2'd2)))))}};
  localparam signed [3:0] p9 = (({2{(2'd2)}}+{4{(2'd1)}})==={1{{3{{1{(2'sd1)}}}}}});
  localparam signed [4:0] p10 = (((5'd27)<(3'sd1))^~((-2'sd1)>(2'd1)));
  localparam signed [5:0] p11 = (!((5'd3)<<(4'sd6)));
  localparam [3:0] p12 = (!({(~^(-4'sd2)),((4'd3)?(3'd4):(2'sd1))}==={{3{(5'd0)}}}));
  localparam [4:0] p13 = (~(~(^(~&(|((-5'sd6)|(-3'sd1)))))));
  localparam [5:0] p14 = ((2'd2)^~(6'd2 * (3'd6)));
  localparam signed [3:0] p15 = (~&(-3'sd2));
  localparam signed [4:0] p16 = (-5'sd6);
  localparam signed [5:0] p17 = (({4{(3'd6)}}-(^(3'd7)))<(((-5'sd2)==(-5'sd0))>>>((3'd0)>(-4'sd4))));

  assign y0 = $signed($unsigned((($signed($signed($unsigned($unsigned($unsigned($unsigned($unsigned((p0))))))))))));
  assign y1 = $unsigned({3{{4{p16}}}});
  assign y2 = (4'd2 * (p8<p8));
  assign y3 = {3{(a1-p12)}};
  assign y4 = ($signed((p14?p10:p12))?(5'd22):$unsigned((p10!=b0)));
  assign y5 = ({{(b5|b5)}}>=((~a0)==(b5+b4)));
  assign y6 = ({(&({p15,p10,p2}<=(|(-5'sd7))))}<<<(((p8)>>(~^p17))<=(~|$signed((!p13)))));
  assign y7 = (-3'sd0);
  assign y8 = {(+(~&(+{p16,a0,a4}))),((~|{1{p2}})>>(~|(-3'sd3)))};
  assign y9 = (b1>=b5);
  assign y10 = $unsigned($signed((|$signed((+($signed($signed((~&((~^a1)>(|b1)))))))))));
  assign y11 = ({a0,p5}<=(a3|p3));
  assign y12 = {4{(!p2)}};
  assign y13 = (((6'd2 * b0)<<<(p3^~p15))^((p3!=p10)%a2));
  assign y14 = (p2+p7);
  assign y15 = (^(4'd11));
  assign y16 = (|(~(~&(~^(&p6)))));
  assign y17 = ((-(3'd4))?(p15?b3:p8):((&b4)+{3{b4}}));
endmodule
