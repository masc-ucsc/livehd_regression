module expression_00856(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(-4'sd3)}};
  localparam [4:0] p1 = (~|(^{(((2'd2)?(-3'sd1):(4'd6))!=((-5'sd2)?(5'd13):(-5'sd11))),({(3'd7),(-2'sd0)}?(-(3'sd1)):(-(5'sd9)))}));
  localparam [5:0] p2 = {3{(2'd0)}};
  localparam signed [3:0] p3 = ((2'd3)<<(-3'sd1));
  localparam signed [4:0] p4 = {(((4'd1)>(2'd1))>>((3'd4)<(2'd0))),{((-3'sd2)<<(3'd5))}};
  localparam signed [5:0] p5 = (&(-((2'd3)&(-2'sd0))));
  localparam [3:0] p6 = {{{{3{((4'sd2)?(3'd3):(5'sd7))}}}},({(5'd9),(-4'sd7),(5'd18)}?{4{(3'd6)}}:{2{(5'sd12)}})};
  localparam [4:0] p7 = (((-4'sd5)<<(4'd10))|{4{(3'd7)}});
  localparam [5:0] p8 = (~^(((2'd0)<<<(2'sd0))||(!(~|(3'd5)))));
  localparam signed [3:0] p9 = {1{(5'sd14)}};
  localparam signed [4:0] p10 = (&{1{((2'd1)^(-3'sd2))}});
  localparam signed [5:0] p11 = ((-4'sd6)>(4'd4));
  localparam [3:0] p12 = {((+(2'sd0))<=(!(-2'sd1))),((~(-5'sd1))^(~^(3'd0))),{{(5'sd0),(-2'sd1),(4'd3)},{(3'd5)}}};
  localparam [4:0] p13 = (((4'd4)^(2'sd0))===((5'd7)>>>(4'sd6)));
  localparam [5:0] p14 = (((((5'd19)^(3'd2))===((5'sd11)&(2'sd0)))>>(((2'sd1)==(2'd2))===((4'd9)>>>(-3'sd1))))>(((-2'sd1)|(4'd4))/(-3'sd0)));
  localparam signed [3:0] p15 = (5'd19);
  localparam signed [4:0] p16 = ((~(~&(-5'sd12)))!==((3'sd3)|(5'd3)));
  localparam signed [5:0] p17 = (&(5'sd15));

  assign y0 = (((a1?p3:p5)?((5'd2 * b0)):(p5?b5:a5))^~$unsigned(((b4?b4:b2)?(b2===b0):((p1?p14:a1)))));
  assign y1 = ({3{p8}}?{2{(p5==p4)}}:(p7?p4:p17));
  assign y2 = (|(-2'sd1));
  assign y3 = (((p10<p5)>=(p8^~b1))=={4{{2{p11}}}});
  assign y4 = (p3?b3:p6);
  assign y5 = {{(p10&a5),{b3,p14,p14}},((~|{a4})>=(p9>=p7))};
  assign y6 = (b1?b2:b3);
  assign y7 = (((a1-b1)?$signed(a4):(a2?a4:p10))?$unsigned(((b5)<(a5^b5))):$unsigned(({3{p0}}<<<(b3^~p8))));
  assign y8 = (((-3'sd1)!=={2{(b0>>a2)}})===({(2'sd0),$signed(a5),{b5,a2,b3}}!=((b0<<<b2)?{1{b5}}:{b1,b1,a0})));
  assign y9 = ({(-(^(p15<=a0)))}!={(p4?p15:p12),(a1&&b5),(b0?p8:a3)});
  assign y10 = {1{{2{(~(~^{1{{2{b0}}}}))}}}};
  assign y11 = (({b5,b5}+(a3))!=={(b1<<b4),(a5||a3),{a1}});
  assign y12 = {4{({3{a5}})}};
  assign y13 = ((-5'sd14)?((p17?p3:p15)?(5'd15):(p8-p2)):{(6'd2 * p1),(p5?p10:p16)});
  assign y14 = (~(~|{(~(&(^(p17|p11)))),(-(~|(&(4'd2 * p7)))),(6'd2 * {p1,p6})}));
  assign y15 = {{(b5>>>p12),{p17}},((4'sd7)^(4'd4))};
  assign y16 = (((a1?p16:a1)?(5'd9):$unsigned(b3))?((2'd1)?(-a4):(4'sd7)):(!(3'd6)));
  assign y17 = ((-4'sd2)<(p13/p1));
endmodule
