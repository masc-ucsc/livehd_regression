module expression_00545(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(-2'sd1),(2'd1)},{2{(3'd1)}},(~(~&(2'd0)))};
  localparam [4:0] p1 = ({((5'd21)|(-2'sd1)),((3'd6)==(3'sd1)),(-(3'd0))}&(~^({(4'd9),(-4'sd6)}^((3'sd1)<(3'd6)))));
  localparam [5:0] p2 = (3'd3);
  localparam signed [3:0] p3 = (((5'd20)?(4'd7):(-4'sd6))^~{(3'd7),(2'sd0)});
  localparam signed [4:0] p4 = (((4'sd0)?(5'd31):(4'd15))?((-4'sd3)==(3'sd2)):((5'd19)===(5'sd12)));
  localparam signed [5:0] p5 = {((2'd3)&&(4'd3)),(4'd2 * (2'd0)),((-2'sd0)&(-4'sd4))};
  localparam [3:0] p6 = (3'sd3);
  localparam [4:0] p7 = ((~^(3'd2))^(2'd2));
  localparam [5:0] p8 = (((4'd2 * (5'd21))+((-5'sd14)>>>(5'd19)))>>>(5'd23));
  localparam signed [3:0] p9 = (((&((4'd3)<(3'd7)))!=((-3'sd0)<=(3'd3)))<=((~^((-5'sd5)===(5'd2)))>=((3'd5)?(3'd3):(4'sd5))));
  localparam signed [4:0] p10 = ((!((-3'sd3)*(-5'sd4)))?((~^(-3'sd2))>(~(-2'sd1))):(~&((-4'sd1)+(3'd7))));
  localparam signed [5:0] p11 = {{(4'd10)}};
  localparam [3:0] p12 = {(-3'sd3)};
  localparam [4:0] p13 = (|((5'd24)+(3'd2)));
  localparam [5:0] p14 = (((2'd3)|(2'd0))?(3'd3):((5'd18)*(5'd3)));
  localparam signed [3:0] p15 = ((4'd7)^~(2'd3));
  localparam signed [4:0] p16 = ((((3'd3)>(5'd30))<{(5'sd1),(4'sd5)})^({(-3'sd0),(2'd3)}&(5'sd8)));
  localparam signed [5:0] p17 = (+((+(-((2'sd0)<<(-4'sd7))))>>(!(~&(^((-5'sd11)!==(-5'sd11)))))));

  assign y0 = (2'd3);
  assign y1 = {p11};
  assign y2 = (p2?p16:a2);
  assign y3 = (({p16,p0,b4}&&(p0?p8:p0))?(~(p8&p11)):((p13?p16:p3)&&{p1,a0}));
  assign y4 = {1{(a3?a1:p12)}};
  assign y5 = $signed((~^(|{(6'd2 * {p1,p13,p1})})));
  assign y6 = $signed(((5'sd12)>=$unsigned(((3'd6)))));
  assign y7 = ($signed({1{(b4|a5)}}));
  assign y8 = (~(!(2'd1)));
  assign y9 = (!(~|((!{1{((a5?a2:b3))}})?{4{(a0^~a3)}}:({p17,a5}?(p9?b5:b3):{a4}))));
  assign y10 = ((p4?p15:p12)&&(p10&p3));
  assign y11 = $unsigned($signed((((b5?b3:a0)?(p3<<<b4):$signed(a2))?(-({3{a2}})):((p16<<<a3)-{3{p1}}))));
  assign y12 = {3{a4}};
  assign y13 = {1{(-5'sd6)}};
  assign y14 = ((p14+p11)^(~^(p0<=p4)));
  assign y15 = ((b2<=a3)*(5'd23));
  assign y16 = (3'd3);
  assign y17 = ($unsigned((4'd2 * {p7,p8,p1}))<((p11>p12)?(~|(p0<p15)):{$signed(p9)}));
endmodule
