module expression_00269(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(|(2'sd0)));
  localparam [4:0] p1 = (~|(~|(~^{3{{4{(4'sd4)}}}})));
  localparam [5:0] p2 = ((((2'd3)>>>(2'd1))?(~^(3'd3)):(~|(2'sd0)))?(((3'sd1)===(5'd21))?((4'd2)>>(5'd12)):((-5'sd10)?(3'd5):(-5'sd4))):((|(-4'sd2))<=((-4'sd3)^~(2'd0))));
  localparam signed [3:0] p3 = (~|(~&(((&(3'sd1))^((2'd2)?(-4'sd0):(5'd15)))>(3'd5))));
  localparam signed [4:0] p4 = (((-2'sd1)-(-4'sd5))?((5'd7)<<<(2'd2)):((4'd11)%(-3'sd1)));
  localparam signed [5:0] p5 = (4'sd6);
  localparam [3:0] p6 = (^(~&{(4'd5)}));
  localparam [4:0] p7 = (({1{(5'd17)}}>=(-5'sd6))<=(((4'd12)>>(2'sd1))|(5'd22)));
  localparam [5:0] p8 = {4{{{{(4'd3),(2'd1),(-5'sd1)}}}}};
  localparam signed [3:0] p9 = ((((5'd12)<(3'sd1))+((3'd5)&(-3'sd2)))<<<({(2'd1),(2'sd0)}^((5'sd12)===(5'd18))));
  localparam signed [4:0] p10 = (~&{1{{2{{3{((2'd3)+(-2'sd1))}}}}}});
  localparam signed [5:0] p11 = (5'd2 * {(4'd7),(2'd2)});
  localparam [3:0] p12 = ((+{{(+(+(~(5'sd4))))}})&&{1{({(4'd6),(3'd3),(-4'sd3)}>=(|((-2'sd1)&&(5'd26))))}});
  localparam [4:0] p13 = ((+(+((4'd11)&(-2'sd1))))&&(~(+(~(-4'sd4)))));
  localparam [5:0] p14 = (3'sd0);
  localparam signed [3:0] p15 = ((~(5'd2 * (~&(5'd27))))<((~^(-3'sd1))|((3'd7)<=(3'd7))));
  localparam signed [4:0] p16 = {1{{3{(5'd2 * (^(2'd1)))}}}};
  localparam signed [5:0] p17 = (((|(~|(5'sd9)))!=((2'd0)!=(-2'sd0)))<((~&((2'd0)===(5'sd1)))<((-3'sd3)*(2'd1))));

  assign y0 = (((2'd2)?(p9&a0):(p2?p3:b3))==(((p7>=p9)&(6'd2 * p2))-((b3>>b4)===(b0&b5))));
  assign y1 = ((((p1*a5)-(5'd26))+(~^(p5-b3)))<<<(&((4'd12)>((p13^p9)>>>(~|p2)))));
  assign y2 = (~^{$unsigned({b5,a0,b2}),{4{p10}}});
  assign y3 = (2'd0);
  assign y4 = (~^(~&p9));
  assign y5 = (~|(((~&b1)|$unsigned(p10))-(2'sd0)));
  assign y6 = ((b4!=a2));
  assign y7 = (((p3&b0)?(-2'sd1):$unsigned(a4))>>(5'd15));
  assign y8 = (3'd5);
  assign y9 = (p5>b0);
  assign y10 = (({4{a5}}?(b5?a0:p8):(p9?b4:b3))?((p4>p17)+{2{b1}}):(5'd2 * (b1+p12)));
  assign y11 = ((5'd4));
  assign y12 = ((p9?p1:p8)*(b1!=b3));
  assign y13 = ({$signed((a5?b2:p5)),(a2>>a0)}?((p11-b4)<={b1,p7,p6}):({p17}?(b2<=p7):(b2==b5)));
  assign y14 = $signed(((-3'sd0)<<($unsigned((p2<<p13))<(p12&&p6))));
  assign y15 = ((~^(~&((|p16)||(p16?a5:p9))))<<<{2{(p2?a0:p2)}});
  assign y16 = {(~|((-(p15&&b1))|({b0,b3,a5}))),($signed((b0<<a1))-(~|{b3,b1}))};
  assign y17 = ((p1?p6:b3)?({a4,b1,b1}!=={a0,a4}):{p13,p10,b0});
endmodule
