module expression_00549(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&{(-3'sd1)});
  localparam [4:0] p1 = {3{(5'd0)}};
  localparam [5:0] p2 = ({{(2'sd0),(-4'sd4),(3'sd0)},((2'd1)>>>(2'd1)),(-3'sd2)}=={(4'd6),(~&(3'sd1))});
  localparam signed [3:0] p3 = ((((4'sd2)!=(-4'sd0))<<<(-3'sd0))>>(3'd4));
  localparam signed [4:0] p4 = ((2'd0)==((4'd14)%(3'sd0)));
  localparam signed [5:0] p5 = (~|(((4'd5)==(-5'sd12))?((5'd23)?(3'd6):(3'd7)):{(-5'sd0)}));
  localparam [3:0] p6 = {({(-5'sd13)}+((-3'sd3)<<(3'd7))),{((5'sd9)-(4'd7)),{(2'sd1)}}};
  localparam [4:0] p7 = (&{(!({(5'd1),(2'd0),(3'sd2)}&&{(4'd0),(3'sd1)})),(|(~&(~(~&{(3'sd0),(2'd0)}))))});
  localparam [5:0] p8 = ((-4'sd5)>>>(-4'sd1));
  localparam signed [3:0] p9 = (~^(((4'd7)||(-3'sd0))<=(~&((5'd23)?(-3'sd1):(5'sd2)))));
  localparam signed [4:0] p10 = {3{(5'sd15)}};
  localparam signed [5:0] p11 = ((~(-3'sd0))<{(5'd0),(2'd3)});
  localparam [3:0] p12 = {((5'sd2)!==(-5'sd4)),((3'sd3)^~(4'd14))};
  localparam [4:0] p13 = {3{((-3'sd2)==(4'd3))}};
  localparam [5:0] p14 = (&(!{{(-4'sd7),(3'd0)}}));
  localparam signed [3:0] p15 = {2{(~^(3'd1))}};
  localparam signed [4:0] p16 = ((3'd5)<={(~&((3'd4)|(3'd6)))});
  localparam signed [5:0] p17 = ({2{(5'd7)}}>>>((4'd0)<<(5'd23)));

  assign y0 = $unsigned((!(~^$signed((~&(4'd3))))));
  assign y1 = ((p13*p1)^(p17^p15));
  assign y2 = ({2{(a0|a5)}}!==(~^{2{{b2,b3,a2}}}));
  assign y3 = ((b3&b0)==(b1&b0));
  assign y4 = $unsigned((5'd2 * (b0&&p8)));
  assign y5 = (5'd18);
  assign y6 = {{a0,b0,a4},{b1,b0,p7},(b4<a1)};
  assign y7 = (($signed(p11)-$signed(a1))?{2{(a2?p15:b0)}}:(-$signed($unsigned(a2))));
  assign y8 = ({p6,b4,a2}?{1{(b4?b0:b3)}}:(p2?a2:b1));
  assign y9 = ((p11>>p6)==(a4>>>p3));
  assign y10 = {a3,a3};
  assign y11 = (~|(a5<<b1));
  assign y12 = {2{(-(~^(((a1?a0:b3)===$unsigned((-a3))))))}};
  assign y13 = ((2'd2)!==(a1?b3:a1));
  assign y14 = {4{p14}};
  assign y15 = (((b4<<<b0)?{2{a3}}:(p14?p6:a4))?((a5&&a1)?(b3<=b5):(b1+p16)):((b3^b3)?{2{b0}}:(b1-b3)));
  assign y16 = {3{((p11<p1)&&(p13|p16))}};
  assign y17 = (-(+{a3}));
endmodule
