module expression_00953(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(^((5'sd5)>>>(2'd2))));
  localparam [4:0] p1 = ((6'd2 * ((5'd6)<<<(3'd6)))?({(4'sd6),(-2'sd1)}>={4{(2'd0)}}):{(-2'sd0),(3'sd1),(5'sd6)});
  localparam [5:0] p2 = {(-4'sd3),(2'd2),(5'd0)};
  localparam signed [3:0] p3 = {{(3'd4),(4'd4)}};
  localparam signed [4:0] p4 = ({2{(!((4'sd5)&(-2'sd0)))}}^~(5'd20));
  localparam signed [5:0] p5 = {{2{((4'd9)?(-4'sd5):(3'd1))}},(5'd2 * {{4{(4'd9)}}})};
  localparam [3:0] p6 = {2{(5'd14)}};
  localparam [4:0] p7 = (((5'd26)<<(2'd2))-((5'd16)&&(5'd30)));
  localparam [5:0] p8 = (|(4'd2 * (2'd1)));
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = (~|(({((2'sd1)?(-2'sd0):(-4'sd4))}||(~^((3'd2)&&(-2'sd1))))-{(&((3'd5)?(5'sd3):(2'd3))),((4'sd7)||(2'd0))}));
  localparam signed [5:0] p11 = {2{((5'sd12)?(4'd5):(-4'sd5))}};
  localparam [3:0] p12 = ({(2'd1),(3'd5)}?((5'd4)?(4'd8):(4'sd4)):((-5'sd12)>>(5'd25)));
  localparam [4:0] p13 = (|(~^(~|((&((3'sd2)^~(-5'sd6)))|(&(~&(-4'sd3)))))));
  localparam [5:0] p14 = {(3'sd0)};
  localparam signed [3:0] p15 = {{(3'd2),(3'd2),(4'd12)},{(4'sd1),(5'd12),(3'sd3)},{(4'd6),(4'sd6),(5'sd8)}};
  localparam signed [4:0] p16 = (~^{1{((((-4'sd6)<=(5'd0))?(-(4'd15)):(+(2'd1)))>({3{(-5'sd13)}}^~((5'd6)<=(2'd2))))}});
  localparam signed [5:0] p17 = {(5'd17),(3'd7)};

  assign y0 = {($unsigned((p6-p6))<<(b4^b4)),((p5?p9:p3)^(p13>p7)),$unsigned(((p1<<<p6)!=(p5?p12:p8)))};
  assign y1 = (+((^((b2)?$unsigned(p12):(b1)))?$unsigned(((p1?p6:b3)|(p8?p2:b0))):(&((|a1)>=(a2^p0)))));
  assign y2 = (4'sd0);
  assign y3 = (-({2{{(a1?p2:p10),$signed(b3),(p15^~a3)}}}));
  assign y4 = (a4?p7:b3);
  assign y5 = {{4{{p6,p12}}},{2{(~(|p11))}},{4{(b2+p16)}}};
  assign y6 = (~|((a2?a1:p2)<<(b0<<<a4)));
  assign y7 = (5'd14);
  assign y8 = (!{({{4{(p12<=a1)}}}-((~(-3'sd2))>>>{p5,p12,b3}))});
  assign y9 = {(a5?a2:b0),(b4?b3:b4)};
  assign y10 = {((p8?p13:p4)+(p2?a5:p1)),((b2+p7)^~(p13?p9:p6)),({p7,p2}?{1{p8}}:(b4>=p7))};
  assign y11 = ((4'sd3)===(-4'sd4));
  assign y12 = {1{(-2'sd1)}};
  assign y13 = (~^((~|(^p0))/p7));
  assign y14 = (!{4{$signed($unsigned(p1))}});
  assign y15 = (p2?b4:a0);
  assign y16 = (((b1?b5:a2)<=(b1?a2:b5))?((a5?b3:p10)||(p17?a2:a4)):((p14-a0)?(a1?b4:p9):{2{p9}}));
  assign y17 = ({(&{a5}),(|(~&a2)),(b4>>a4)}==={3{(+(2'd2))}});
endmodule
