module expression_00914(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(3'd0));
  localparam [4:0] p1 = (-(~|(~|(({2{(-2'sd1)}}|((5'd22)^~(2'sd1)))<{1{((5'sd1)+(4'd4))}}))));
  localparam [5:0] p2 = {{{4{{(4'd6)}}},{{2{{(5'sd4),(5'd1),(4'd11)}}}}}};
  localparam signed [3:0] p3 = (~&((4'd2 * (2'd2))||((4'sd6)+(2'd1))));
  localparam signed [4:0] p4 = (((5'sd3)?(4'd8):(-2'sd0))?((-5'sd4)==(2'sd0)):((-2'sd0)+(3'd7)));
  localparam signed [5:0] p5 = (((5'd9)^~(2'sd0))!==(^(3'd3)));
  localparam [3:0] p6 = {1{({2{(2'd2)}}-(~{(4'sd6),(4'sd7),(-3'sd2)}))}};
  localparam [4:0] p7 = {4{((-2'sd1)^~(5'd7))}};
  localparam [5:0] p8 = {(5'd7)};
  localparam signed [3:0] p9 = (((3'd3)-(-3'sd0))+(~&(|(3'd4))));
  localparam signed [4:0] p10 = (-(~|(^(~&(~|(4'd1))))));
  localparam signed [5:0] p11 = ((3'd5)?((5'd21)?((5'sd4)?(4'd1):(4'd11)):((4'sd3)?(4'sd1):(4'd13))):(-2'sd0));
  localparam [3:0] p12 = ({2{(2'd2)}}<<<((3'd3)^~(2'd2)));
  localparam [4:0] p13 = ((((2'd2)<(5'd16))|((3'd1)^~(3'd0)))<<(3'sd3));
  localparam [5:0] p14 = ({1{(^{(3'd3),(4'd15),(4'd3)})}}?{(2'd1),((-3'sd1)?(2'sd1):(2'sd0))}:(~{2{(4'd6)}}));
  localparam signed [3:0] p15 = (3'sd3);
  localparam signed [4:0] p16 = (5'sd3);
  localparam signed [5:0] p17 = ({2{(4'd12)}}|((-3'sd3)!=(2'd3)));

  assign y0 = ({2{{4{p15}}}}&((~|(+(p16|p9)))&(|{4{p10}})));
  assign y1 = (|$signed((($signed((p11?a5:a5))^((~|p17)))^~(5'd2 * (~&$unsigned(a2))))));
  assign y2 = ({1{b5}}?(b4?b3:b0):(b5^b1));
  assign y3 = (~&{4{(3'd2)}});
  assign y4 = (-5'sd14);
  assign y5 = {(+(|({1{$unsigned(((a5)!==(!b1)))}}&$unsigned(((5'd22)^~(-4'sd7))))))};
  assign y6 = $signed(({4{p1}}-(((p0)&$unsigned(p14)))));
  assign y7 = ((((a4!=a3)!==(a0===b4))||(2'd1))|(({a4}===(a4||b1))^((p16>>>b3)<<<(p4+a4))));
  assign y8 = (b1?b0:b2);
  assign y9 = (+(({1{(a3>b2)}}>=(+(b3!==a1)))?(~$signed({{b0},{p14,b2},(a3+b3)})):((p7<=b3)?(+p12):(~b5))));
  assign y10 = ((a2>a2)>>(a3!==b0));
  assign y11 = ((5'd2 * a0)<<{3{a4}});
  assign y12 = $unsigned((5'sd2));
  assign y13 = (&(&{(~|(&(p4<<<p6))),(~(p5?p9:p13)),(p10?p17:p8)}));
  assign y14 = (4'd14);
  assign y15 = (|{{b2},(b5<p0),{4{p3}}});
  assign y16 = ($unsigned((~&p11))>={2{p10}});
  assign y17 = $unsigned(($signed((~&b5))*(a5?p9:b0)));
endmodule
