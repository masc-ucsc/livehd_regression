module expression_00578(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd5)-(5'd8))?((3'd6)?(3'd2):(3'd1)):{1{(2'd2)}});
  localparam [4:0] p1 = ((((-3'sd0)-(5'd7))===((-4'sd0)>>>(4'sd4)))^~(((-4'sd7)?(-5'sd2):(-3'sd3))<((4'd7)===(2'd0))));
  localparam [5:0] p2 = ((((4'd15)?(5'sd9):(4'sd0))^{{((2'sd0)<=(-5'sd14))}})<<{({(4'd12),(5'd28)}||{1{((4'd6)?(-5'sd14):(5'sd5))}})});
  localparam signed [3:0] p3 = (((-4'sd6)||(5'd0))?{(3'd4)}:(5'd23));
  localparam signed [4:0] p4 = (((3'sd1)===(5'd23))>>>((5'sd7)<<(3'sd3)));
  localparam signed [5:0] p5 = ({((5'sd12)-(-5'sd6)),(4'd2 * (5'd10))}&&{((5'd26)^~((-2'sd0)>>(-4'sd4)))});
  localparam [3:0] p6 = (~^(2'sd1));
  localparam [4:0] p7 = (~&(~{4{(~(5'sd1))}}));
  localparam [5:0] p8 = ((((2'sd1)+(4'd14))||((-3'sd3)-(3'd3)))^({(2'sd0),(4'd11),(-3'sd3)}<=((3'sd2)<(4'd5))));
  localparam signed [3:0] p9 = {2{(~(((3'sd1)|(3'sd1))>={3{(-3'sd3)}}))}};
  localparam signed [4:0] p10 = (4'd4);
  localparam signed [5:0] p11 = (((2'd2)^(-4'sd6))>((-2'sd0)?(5'sd15):(4'd11)));
  localparam [3:0] p12 = (3'sd1);
  localparam [4:0] p13 = {((+(((3'd3)+(-4'sd7))>>((3'd6)^~(3'd3))))<(~&(((-5'sd0)<=(4'd13))?{(5'd27)}:{(4'd0),(-2'sd1)})))};
  localparam [5:0] p14 = ((((5'd25)&(4'sd3))|{1{((3'd4)^(4'sd3))}})|(((-4'sd0)<<(2'd1))?((2'd2)>(5'sd1)):((-3'sd3)?(3'd7):(3'sd3))));
  localparam signed [3:0] p15 = (~|(~^(~|((2'd0)?(5'sd6):(5'd2)))));
  localparam signed [4:0] p16 = ((^(~(2'sd0)))?((2'd2)?(-4'sd4):(5'sd10)):(4'sd0));
  localparam signed [5:0] p17 = (~^(4'sd7));

  assign y0 = (-2'sd0);
  assign y1 = (3'd6);
  assign y2 = $unsigned({4{b2}});
  assign y3 = (~&{3{(~^(~&{3{a3}}))}});
  assign y4 = ((3'd5));
  assign y5 = $signed($signed({4{p4}}));
  assign y6 = (-{{(!(-{p9,p9,a2})),{{{p5},{p7,p8},{a4}}},(~&(-(~|{p12,p11,p14})))}});
  assign y7 = (5'd28);
  assign y8 = ((({4{a0}}||(a4?b1:a1))^(a1?p8:b0))+(((a1<<a3))>=((b4||a2)^~(a0?b0:a2))));
  assign y9 = {4{{2{p17}}}};
  assign y10 = ((5'd2 * b0)^$unsigned(p7));
  assign y11 = {{{({b5,b1,a3}!==(a0<=b3)),{{b5},(a5===b4)}},({(2'd0),{b5,a4,b5}}-$unsigned((5'd0)))}};
  assign y12 = (((~|b1)>>>(p8%p15))^~(-4'sd5));
  assign y13 = ($signed(p11)?(a0?p14:p0):(5'd0));
  assign y14 = (5'sd14);
  assign y15 = ((~((~^p6)>>(b5&&p9)))&&(2'd2));
  assign y16 = {1{(({4{b2}}=={2{a2}})+{1{{2{(a1?a3:a0)}}}})}};
  assign y17 = ((-3'sd0)>=(~^(!(~(^(~|(2'd2)))))));
endmodule
