module expression_00326(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd6)?((5'sd15)?(-4'sd4):(3'sd3)):(2'd3));
  localparam [4:0] p1 = (((~(~^(5'd14)))>{((4'd0)+(5'd24))})^~(!(~&{((3'sd3)>>>(-2'sd0))})));
  localparam [5:0] p2 = {(2'sd0),{{(-5'sd6),(4'sd7)}},{(4'sd5)}};
  localparam signed [3:0] p3 = (-4'sd2);
  localparam signed [4:0] p4 = ({(3'd4),(5'd7)}?(~^(2'sd1)):(6'd2 * (5'd25)));
  localparam signed [5:0] p5 = (({3{(5'sd3)}}>((4'sd1)-(2'sd0)))>={4{(2'd0)}});
  localparam [3:0] p6 = (~|({(2'd2),(2'd2)}<<<((~((3'sd2)||(5'sd8)))===(~|(&(2'd1))))));
  localparam [4:0] p7 = (~&((|{4{(-(2'd3))}})&&{3{{(3'd3)}}}));
  localparam [5:0] p8 = ((!(((4'sd2)-(-4'sd7))^((2'sd0)?(2'd3):(4'd2))))?(-5'sd10):((-(-5'sd12))-(-3'sd0)));
  localparam signed [3:0] p9 = ((~|(((4'd5)<<(-2'sd1))<=(^(~&(2'sd0)))))<<({2{{(3'd7),(5'd9),(2'd2)}}}=={(3'd5),(-5'sd12),(4'd2)}));
  localparam signed [4:0] p10 = ((((2'sd1)-(2'sd0))||((-5'sd6)||(3'sd2)))&&{3{(-3'sd3)}});
  localparam signed [5:0] p11 = {(((5'sd15)<<(3'sd0))^~((3'd6)?(4'd4):(4'sd1))),{((3'd1)>>(4'd0)),((5'd28)&&(3'd6))}};
  localparam [3:0] p12 = {4{((-2'sd0)<{(4'sd3)})}};
  localparam [4:0] p13 = {4{{2{(2'd0)}}}};
  localparam [5:0] p14 = (((-3'sd1)?(4'sd4):(-3'sd2))?((3'sd3)<<(2'd1)):((3'd4)==(4'sd7)));
  localparam signed [3:0] p15 = (((4'd0)==(2'sd1))?(((-3'sd2)===(3'd4))<((2'd2)?(-4'sd4):(-2'sd1))):(((5'd0)?(3'sd2):(5'd1))===((2'd0)||(-5'sd4))));
  localparam signed [4:0] p16 = {(+(2'sd0)),((3'sd0)?(5'd1):(4'sd3)),(|(5'd13))};
  localparam signed [5:0] p17 = {((3'sd1)?(3'd1):(4'd8))};

  assign y0 = {2{(3'd1)}};
  assign y1 = ($unsigned(a2)-(4'd2 * p0));
  assign y2 = $unsigned((((a5!=b5)<<<(b4!==a0))^(!{4{(-b4)}})));
  assign y3 = (!(~{b1,b2}));
  assign y4 = (($signed((p1&&p2))&(p16?p17:p3))||(-4'sd0));
  assign y5 = {4{{4{p11}}}};
  assign y6 = ({(a4?b4:a1),(b1||a3),(b3!==a5)}|((b2!=a5)<<{b2,a1,b4}));
  assign y7 = (((~|(b3<<b5))&&$unsigned((+(b2/a4))))<(~|(3'd2)));
  assign y8 = (3'd0);
  assign y9 = ((2'sd0)<=(({3{b3}}===(a3&&a3))>(~|(~&$signed(p10)))));
  assign y10 = $signed($unsigned(p2));
  assign y11 = $signed((5'd16));
  assign y12 = ({$signed({a5,b2,a3}),$signed($unsigned(a1))});
  assign y13 = {1{({p2}<<(~|p10))}};
  assign y14 = (|(^((&(b0-p0))?(b4?p6:p10):(b5?p11:b0))));
  assign y15 = {1{({1{p16}}?(b0^b0):(a1?b1:b2))}};
  assign y16 = {4{((a2>a2)>>(~|a2))}};
  assign y17 = ($unsigned({b2})!==(-{b5,a1,b4}));
endmodule
