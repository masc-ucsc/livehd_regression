module expression_00649(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(^(5'd2 * (~|(4'd5)))));
  localparam [4:0] p1 = ((2'd3)^({(2'd0),(4'sd4),(-5'sd7)}|((5'd14)>=(3'd2))));
  localparam [5:0] p2 = (-3'sd3);
  localparam signed [3:0] p3 = (((6'd2 * (5'd17))?((2'd1)?(2'd3):(2'd3)):((2'd2)%(4'sd4)))-(((4'd6)<<(4'sd4))-((2'sd0)==(-5'sd6))));
  localparam signed [4:0] p4 = (5'd2 * ((3'd6)-(5'd18)));
  localparam signed [5:0] p5 = (^({3{(2'd0)}}?{4{(4'd13)}}:{4{(3'd3)}}));
  localparam [3:0] p6 = (^(3'd2));
  localparam [4:0] p7 = ({(+((-2'sd0)>=(2'd0))),{(5'sd1),(-3'sd0),(3'd5)}}|({(2'sd0),(4'sd7)}&((2'd0)<(3'sd0))));
  localparam [5:0] p8 = ({4{(-3'sd3)}}?(3'd3):{(-3'sd2),(-4'sd2),(-5'sd1)});
  localparam signed [3:0] p9 = ((((-3'sd2)==(4'd6))?((-5'sd3)?(5'd0):(2'sd0)):((5'sd14)&&(4'sd2)))?(((-3'sd2)|(2'd1))<<((4'd6)?(-2'sd0):(3'd4))):((5'd2 * (5'd2))<<<((5'd17)?(4'd1):(5'sd2))));
  localparam signed [4:0] p10 = (!(~|{{2{{((2'sd1)>>>(2'd1))}}}}));
  localparam signed [5:0] p11 = ((3'sd0)==(3'd7));
  localparam [3:0] p12 = ({(2'd3),((2'd3)&&(3'd3)),(2'd3)}!==(~(~&(|(((5'd30)>(5'd27))+(~^(3'd3)))))));
  localparam [4:0] p13 = ((((-3'sd2)?(5'sd9):(5'sd2))||(5'sd6))>((-4'sd5)<<(3'd1)));
  localparam [5:0] p14 = ({4{((5'sd1)<(3'sd0))}}-{2{((4'd4)>(5'd30))}});
  localparam signed [3:0] p15 = ({2{{(3'd7),(3'd3),(4'd11)}}}+{4{(2'd1)}});
  localparam signed [4:0] p16 = (|(&(4'sd5)));
  localparam signed [5:0] p17 = ((((4'sd1)==(3'sd2))^((4'd9)<=(4'd8)))>=(((2'd1)&(4'd10))>>>((3'd5)||(2'sd0))));

  assign y0 = ({(&(-2'sd1))}<<<(2'd1));
  assign y1 = {((4'sd0)^(+(^((p5?p5:p17)<<(p3?p3:p14)))))};
  assign y2 = (-(&{(&$signed({{p14,a2}})),(~{(^a2),$unsigned(a0),(a1)})}));
  assign y3 = {4{a5}};
  assign y4 = ((a3?p16:b5)<<(4'd7));
  assign y5 = (({a5,a3}&(a3||a4))!==(5'd2 * {b2}));
  assign y6 = $unsigned(({2{a1}}>>{p12,b0,b2}));
  assign y7 = (!(-{2{((~(a3))?(a5&&a3):(p0?b4:a4))}}));
  assign y8 = {2{(~|(^(^{2{{2{b1}}}})))}};
  assign y9 = $signed(($unsigned({2{b3}})));
  assign y10 = (((&(p15!=a0))>(-3'sd1))>$signed((2'd3)));
  assign y11 = {{{p15,b3,p15},(b0!==a2),(b0&&p10)},$signed(($signed({(a0>=b0)})!=={b0,a3,b2}))};
  assign y12 = {((a4^~b1)|(!a3)),({a1,a0,b0}==(-b0))};
  assign y13 = ((p12-p9)>>(p7^~a5));
  assign y14 = ((p14>>p9)|(5'd2 * p8));
  assign y15 = $unsigned((!b3));
  assign y16 = {b3,b5,a0};
  assign y17 = {1{{1{{4{(!(&{3{p15}}))}}}}}};
endmodule
