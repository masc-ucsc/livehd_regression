module expression_00055(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {({(3'sd3),(-5'sd0)}>>>((4'd4)?(-3'sd1):(5'd13))),{{{(-2'sd0),(2'sd0)},((3'd4)&&(5'd30)),{(3'd4),(4'd9),(2'd0)}}}};
  localparam [4:0] p1 = (((-3'sd0)>>(5'd12))?(~&((2'sd1)===(2'd3))):(~^(~&(4'sd3))));
  localparam [5:0] p2 = (!(~(!(&(~&(^(~&(&(~(|(!(~|(-2'sd0)))))))))))));
  localparam signed [3:0] p3 = (~|(!{1{(+({4{(-5'sd9)}}>((&(3'd3))||{(2'sd1)})))}}));
  localparam signed [4:0] p4 = {3{((~^(5'sd5))||{1{(5'd24)}})}};
  localparam signed [5:0] p5 = (((4'd10)^~(2'd0))&&(~|((5'd31)||(3'sd3))));
  localparam [3:0] p6 = {4{((2'd1)&&(2'd2))}};
  localparam [4:0] p7 = ({(2'd2),(-4'sd7),(5'd30)}?{(2'sd0),(3'd1)}:((3'd1)?(-4'sd0):(2'd0)));
  localparam [5:0] p8 = (((-2'sd1)?(5'sd0):(5'd8))?((5'd18)?(2'sd0):(3'sd0)):((3'd3)?(2'd0):(2'd2)));
  localparam signed [3:0] p9 = ({2{(4'd6)}}>>>((2'sd0)<(4'd1)));
  localparam signed [4:0] p10 = (2'sd0);
  localparam signed [5:0] p11 = (({(-(5'sd11))}?(5'd2 * (4'd9)):((3'd7)<<<(3'd4)))^(((4'd6)==(5'd28))?(~^((3'd4)||(4'd2))):(~|((3'd0)&(3'sd0)))));
  localparam [3:0] p12 = {{{((4'd14)<=((-4'sd7)<=(4'sd6)))},((~|(5'd14))&((-2'sd1)||(3'd5)))}};
  localparam [4:0] p13 = (~^{2{(4'd2 * (~|(~^(4'd3))))}});
  localparam [5:0] p14 = ((5'd12)?(&(4'd12)):((3'd6)-(4'd11)));
  localparam signed [3:0] p15 = {1{({{(5'sd8),(4'sd0),(5'sd0)},((-4'sd1)<<<(-5'sd10)),{4{(2'd2)}}}>>>(6'd2 * ((4'd0)!=(5'd29))))}};
  localparam signed [4:0] p16 = {((^(4'd15))?(+(4'd9)):{(-4'sd4),(5'd26)}),((~^(5'd4))?(~^(-4'sd4)):{(3'sd2),(-3'sd2),(-3'sd2)}),(2'sd0)};
  localparam signed [5:0] p17 = ((-4'sd1)^~(-3'sd1));

  assign y0 = {3{{p2,p2}}};
  assign y1 = {{$unsigned(b1),{a5,b3}},(5'sd15),((5'd31))};
  assign y2 = (-((+(2'sd1))&(b1>=b4)));
  assign y3 = (~^(+((-4'sd2)<<<$unsigned(b2))));
  assign y4 = $unsigned((((~&$signed((~^(!(&p1))))))));
  assign y5 = (|((~(((~&{1{{4{a2}}}})+$unsigned((|(a0||b1))))!==((^(^{3{b5}}))-($unsigned(b5)>>(!b4)))))));
  assign y6 = (((a2?a4:a1)!==(a5-a1))?((p2>>p8)>={(3'sd2)}):({1{p4}}?(-3'sd2):(a3|b1)));
  assign y7 = ((&((b1<p10)))^~((a1?a2:a0)&$unsigned(p11)));
  assign y8 = (6'd2 * (p14?b1:b1));
  assign y9 = (~|(~|(($unsigned((4'd8)))!==(~((3'sd0))))));
  assign y10 = (4'd10);
  assign y11 = (2'd1);
  assign y12 = (4'd12);
  assign y13 = (a4^b5);
  assign y14 = {2{((a4<=b2)<<(p8-p11))}};
  assign y15 = (((b0<=p16)?(a5?a5:a2):(a5==b5))!=((a1?a4:a4)>>(b0-b0)));
  assign y16 = $signed(($unsigned((a0>>p3))^$signed((p10+a5))));
  assign y17 = ({(a1?b1:b4),(~&(p17?b2:a0))}?(~&{(&(4'd2 * a0))}):((a2?b2:p1)?(p15>=a1):(a1?a2:b1)));
endmodule
