module expression_00500(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-2'sd0);
  localparam [4:0] p1 = {{({3{(-2'sd0)}}<=((-4'sd4)+(2'sd1))),{4{(3'd1)}},(((4'd13)?(-4'sd5):(-5'sd11))|{(5'sd6)})}};
  localparam [5:0] p2 = (({3{(2'd2)}}|{4{(-5'sd14)}})<<<{3{(4'd12)}});
  localparam signed [3:0] p3 = ((5'd20)||(5'd17));
  localparam signed [4:0] p4 = {2{(!((4'd4)?(4'd5):(-2'sd1)))}};
  localparam signed [5:0] p5 = (~|(&(-2'sd1)));
  localparam [3:0] p6 = {(~^(3'd6)),((3'd2)?(5'sd4):(-5'sd7))};
  localparam [4:0] p7 = (((4'sd0)==(2'd3))?((-2'sd1)>>>(4'sd0)):((5'sd1)?(5'd15):(3'sd2)));
  localparam [5:0] p8 = (~((3'd4)+((~(4'sd5))^(-3'sd0))));
  localparam signed [3:0] p9 = ((((2'd3)&&(-5'sd8))?{(3'd7),(4'sd6),(-5'sd6)}:((2'd1)-(5'd28)))?(((5'sd2)-(-3'sd2))?(!(2'd3)):{(3'd4),(2'd0)}):(((3'd7)?(-3'sd1):(2'd3))?((-3'sd2)-(3'd0)):(~(2'd3))));
  localparam signed [4:0] p10 = (2'sd0);
  localparam signed [5:0] p11 = ((-5'sd13)||(4'd15));
  localparam [3:0] p12 = {4{(~|(~|(~^(-3'sd3))))}};
  localparam [4:0] p13 = ({(-2'sd0),(5'd18),(3'd6)}-(((-5'sd5)>>>(2'sd0))<<<{(3'd7),(4'sd4)}));
  localparam [5:0] p14 = ((((-3'sd0)===(5'd11))<<((2'sd0)<=(5'd28)))!=={2{((4'd10)^(5'd1))}});
  localparam signed [3:0] p15 = ((4'd2)<<((2'd1)?(4'sd4):(-5'sd9)));
  localparam signed [4:0] p16 = ({4{(-3'sd0)}}<=(^((3'd1)&&(-5'sd2))));
  localparam signed [5:0] p17 = (((5'd26)+(2'd1))<((-5'sd7)^~(3'd2)));

  assign y0 = (^$signed(({3{{2{p7}}}})));
  assign y1 = ({2{b4}}?(p5|a0):{3{p0}});
  assign y2 = ((&(~|p4))<={b1,b2,b4});
  assign y3 = {{a0,a0,p4},(~|(p9?a1:b2)),(!(~&(a0^b3)))};
  assign y4 = {3{{a2,p4}}};
  assign y5 = (3'd1);
  assign y6 = (~&(+(((b4-b0)<(b1^~b4))==={1{((4'd2 * b2)!=={4{a1}})}})));
  assign y7 = (((a5?b0:p1)-((a2?b5:b5)===(!b3)))-((+(p8?a5:b3))?(a4||b3):(p8?a5:b5)));
  assign y8 = {((~|(+(((b5===b5)==(a0+p8))&{$signed((~^{(-(|p6))}))}))))};
  assign y9 = ((!(b0>=b1))-(~&(p12|p6)));
  assign y10 = {4{((|p11)>>>(~|p3))}};
  assign y11 = ((|(p1>p16))<((p4/p4)+(-p13)));
  assign y12 = {((~^{p17,p14})>=$signed({a5,p7}))};
  assign y13 = (3'sd1);
  assign y14 = ((((~|a3)||{2{a0}})===(~((5'd2 * b0)<(~&a4)))));
  assign y15 = ((|p5)==(-p12));
  assign y16 = {(5'd2 * p7),(p8>>>p4),{p16,p16}};
  assign y17 = (!(5'sd13));
endmodule
