module expression_00780(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(2'd3),(4'sd0)}};
  localparam [4:0] p1 = (~&(|(-2'sd1)));
  localparam [5:0] p2 = (((3'sd2)-(4'd2))+((3'sd0)?(3'd6):(3'd3)));
  localparam signed [3:0] p3 = (({(2'd0),(5'sd8)}>>((-4'sd4)+(5'sd13)))!=={((-3'sd2)^~(-3'sd3)),((4'd1)>=(3'sd1)),{(5'd22),(-4'sd7),(-4'sd1)}});
  localparam signed [4:0] p4 = {1{({1{(-4'sd1)}}!=={2{(3'd4)}})}};
  localparam signed [5:0] p5 = (4'd10);
  localparam [3:0] p6 = ((4'd14)?(-4'sd0):(5'd10));
  localparam [4:0] p7 = ((((-4'sd2)>=(5'd14))?((2'd1)&(4'd7)):((2'sd1)?(-2'sd1):(5'd10)))?(((5'sd13)^(2'd3))?((2'd2)?(5'sd4):(2'd0)):((4'd13)==(4'sd7))):(((4'd0)?(-2'sd0):(-2'sd1))&&(+(-2'sd1))));
  localparam [5:0] p8 = (4'sd1);
  localparam signed [3:0] p9 = {1{{3{((2'd3)?(4'sd1):(3'd7))}}}};
  localparam signed [4:0] p10 = (({(4'sd2),(3'd3),(-5'sd9)}|((3'd6)&&(2'sd1)))<{(2'sd1),(-3'sd3),(3'd0)});
  localparam signed [5:0] p11 = (((3'd2)>(5'd26))?((3'd6)<(4'd8)):((-5'sd11)||(4'd7)));
  localparam [3:0] p12 = ((-(!((4'd3)?(4'd5):(5'sd14))))?((~^(-2'sd1))?((3'sd3)&&(5'sd3)):((2'sd0)+(4'd14))):(6'd2 * ((2'd0)?(4'd11):(2'd0))));
  localparam [4:0] p13 = (-((~^(4'sd1))>>((-2'sd1)?(2'd0):(3'd0))));
  localparam [5:0] p14 = {(4'd15)};
  localparam signed [3:0] p15 = (~|(((5'd18)<<<(3'd4))?(^(-3'sd0)):{(-3'sd0),(3'd6)}));
  localparam signed [4:0] p16 = (|({{3{(2'sd1)}},(^(-5'sd13)),(5'd9)}<<<(((3'd1)+(4'd15))<<<{(5'sd0),(5'd31),(4'd9)})));
  localparam signed [5:0] p17 = ((&(4'd13))^~(-3'sd1));

  assign y0 = ((-b0)?(^b4):(p15?a4:b5));
  assign y1 = {4{{3{{a2}}}}};
  assign y2 = ((4'd2 * (p0<=p7))<=({3{p6}}<<{4{p9}}));
  assign y3 = {p4};
  assign y4 = {{2{{p1,p9,p12}}},{4{(a5?p15:b5)}},(+{3{(p11?p1:b4)}})};
  assign y5 = (~&{2{{b3,b2,b3}}});
  assign y6 = {a0};
  assign y7 = {3{{p1,b1,p17}}};
  assign y8 = {$signed(b4),(4'd8)};
  assign y9 = (a0!==b3);
  assign y10 = (((-((a0===b0)>>(|b5)))&((!a4)===(a3<b2)))+(5'sd9));
  assign y11 = (b3>p14);
  assign y12 = (-5'sd10);
  assign y13 = ((p2?b2:b2)?(p13?b2:a0):{{p0,p17,p6},(p6?b1:p5)});
  assign y14 = ({3{{2{a2}}}}!==({3{(~&a3)}}!==((a2>>b3)&&(~^a0))));
  assign y15 = $unsigned((~|((p1<<<p8)&(a4>p1))));
  assign y16 = ({4{b5}}!==(b1!==a1));
  assign y17 = (4'd11);
endmodule
