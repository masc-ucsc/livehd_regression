module expression_00215(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{4{(4'd7)}}}};
  localparam [4:0] p1 = (5'd19);
  localparam [5:0] p2 = ({3{((4'd6)<=(-5'sd2))}}!==(^((~|(-4'sd3))<<((5'sd12)|(-4'sd2)))));
  localparam signed [3:0] p3 = {1{({4{(4'sd1)}}>=(~&(2'd0)))}};
  localparam signed [4:0] p4 = {1{{4{(4'd13)}}}};
  localparam signed [5:0] p5 = (+(~({(&(3'd7)),((3'd0)===(5'd24))}|({3{(2'd2)}}==(3'd1)))));
  localparam [3:0] p6 = (~&{(3'd0),(-2'sd1)});
  localparam [4:0] p7 = (5'sd11);
  localparam [5:0] p8 = (({(2'd3),(5'd16)}?((2'd2)!=(5'd5)):{(5'd19)})<({(5'sd6),(3'd0),(2'sd1)}?(-5'sd15):((4'd12)?(-4'sd6):(-2'sd0))));
  localparam signed [3:0] p9 = {(4'sd4)};
  localparam signed [4:0] p10 = ((((5'd25)!==(5'sd6))^~(^((5'sd9)>>(5'd19))))-((~{1{(5'd20)}})&&(^((-3'sd2)===(5'd15)))));
  localparam signed [5:0] p11 = {(~|(+(~(~^(4'd10))))),{(-(4'sd6)),(~&(3'sd1))}};
  localparam [3:0] p12 = ((~|((^(-3'sd3))!==((3'sd1)===(2'sd0))))+(4'd14));
  localparam [4:0] p13 = {2{(5'd11)}};
  localparam [5:0] p14 = (&{{2{(-2'sd1)}},{1{((2'sd0)^~(-4'sd1))}},{1{((-4'sd4)!=(4'd7))}}});
  localparam signed [3:0] p15 = {(|(~|(~^(~|(2'sd1)))))};
  localparam signed [4:0] p16 = (~&((-(2'd0))>>>(5'd28)));
  localparam signed [5:0] p17 = ((4'd2 * (&((2'd2)||(4'd7))))>(~|({(2'd3),(3'sd1),(-5'sd7)}^(!(5'sd14)))));

  assign y0 = (4'd4);
  assign y1 = (-4'sd1);
  assign y2 = ((2'd0)^(4'd7));
  assign y3 = {p4,p7,p12};
  assign y4 = ((~&(~&{a4,p12}))<<<{{2{p7}},(~^p2),(b1<p16)});
  assign y5 = (a4|a4);
  assign y6 = (-p2);
  assign y7 = (^(+(~(+(|(~^(!((b2>p11)^(!(p13%p15))))))))));
  assign y8 = (&({(p13>>p16),(|a0),(a1^~p12)}>>((b1&&p7)^{p13,p0,a4})));
  assign y9 = {(5'd20),((5'd27)&(p4^~p10)),{(5'sd7),{p14,p2}}};
  assign y10 = ({({p11}<=(p1||p5)),({b1,p0,p4}^~(p4-p4))}|{{(p16>a4),(a4>>p17),(b4+p9)}});
  assign y11 = (~^(&($unsigned($unsigned(a4))>=(a2>>b4))));
  assign y12 = ({1{(~&$signed({1{(({2{b0}}?{a2,a0,p5}:(+p12))?$unsigned($unsigned((p7?p13:b4))):((b0?p14:b4)))}}))}});
  assign y13 = $unsigned({((3'd1)),$unsigned((4'sd4))});
  assign y14 = ((({a1}?{p5,a2,b3}:(b5<a0))|((4'd2 * a0)?{a5}:{a3,b3}))=={({a2,p4}^~(b5<<<a4)),{((a5?b1:p13)<<(b2===a2))}});
  assign y15 = ((^(((p11<<<p1)>>$signed(a3))+(!{2{p4}})))<<{1{((|$signed((((^p16)<<(~&p3))))))}});
  assign y16 = ({a5}?(a2?p0:a4):{4{a3}});
  assign y17 = {3{{1{(b3?b1:a0)}}}};
endmodule
