module expression_00687(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(5'd15)};
  localparam [4:0] p1 = ((((2'd2)?(5'd20):(4'd6))>>((4'd11)-(-3'sd0)))?{((2'sd1)<=(4'd4)),((2'd3)|(-5'sd8)),((4'd12)||(3'd5))}:{4{(5'sd8)}});
  localparam [5:0] p2 = ((&(^(~(~&(4'sd5)))))<<(^(~|((4'd15)==(3'd1)))));
  localparam signed [3:0] p3 = (2'd1);
  localparam signed [4:0] p4 = (-{{{(2'd2),(4'd3)},{(5'd6),(-2'sd0)},{(3'd3),(5'd6),(-5'sd0)}}});
  localparam signed [5:0] p5 = (((-(-3'sd2))?(~&(2'd1)):(~(-2'sd0)))>((^((3'd2)!=(3'd3)))>=((-4'sd2)?(-5'sd4):(5'd7))));
  localparam [3:0] p6 = (2'sd0);
  localparam [4:0] p7 = ((&(!((-(4'd0))&((2'd1)>>>(3'd4)))))&&({{2{(3'd7)}}}|{(3'sd3),(2'd0)}));
  localparam [5:0] p8 = ((((3'd6)?(5'd16):(3'd5))==((-5'sd9)?(5'sd11):(-5'sd11)))?(((2'd1)>(-2'sd1))===((-2'sd1)<<(4'sd0))):(((2'sd0)>>>(5'd6))&((-3'sd0)?(2'sd1):(4'd2))));
  localparam signed [3:0] p9 = (((5'd15)<((-4'sd1)+(3'd1)))|({1{(3'd1)}}?((2'sd1)?(4'd5):(4'd0)):{(3'd3)}));
  localparam signed [4:0] p10 = (((-3'sd0)?(-3'sd2):(3'sd3))?(((-2'sd0)?(-5'sd15):(3'd7))+(~|(2'sd1))):((4'd9)?(5'd2):(3'sd3)));
  localparam signed [5:0] p11 = (~&(~|(~(4'd0))));
  localparam [3:0] p12 = (~&(5'd5));
  localparam [4:0] p13 = {(-4'sd7),(~^(2'd2)),{4{(4'd8)}}};
  localparam [5:0] p14 = ({((3'sd0)^(5'd8))}&&{((3'd3)&&(3'd0)),{(3'sd1)},(4'd2 * (4'd13))});
  localparam signed [3:0] p15 = (!(4'd13));
  localparam signed [4:0] p16 = (3'sd2);
  localparam signed [5:0] p17 = {({(-5'sd13),(2'd1)}||((3'sd2)!=(2'd0))),{(~(5'd26)),(!(-5'sd14))}};

  assign y0 = (!((b0===b4)|{p16,a5}));
  assign y1 = (!(~^(4'd11)));
  assign y2 = (($unsigned((p1-b5))|(b5?p9:a0))^((a0?b1:b2)?$signed((p12==b1)):$unsigned((p4?p6:a1))));
  assign y3 = ((p5?a4:p11)?((p8)/p6):(~(~^(p15^p9))));
  assign y4 = ((a5-b1)?(b1?a2:p16):(-(p1?a5:p13)));
  assign y5 = $unsigned(({{p2,p15,p12},(p10+p6)}||({p12}||(p7^~p11))));
  assign y6 = (4'd2 * p14);
  assign y7 = ({p15,p13}^~(^p3));
  assign y8 = $signed({3{($unsigned(p10)>>(p0))}});
  assign y9 = (^$signed((($unsigned(b5)||(-4'sd4))?(a2?b3:p6):{2{{b0}}})));
  assign y10 = (~^{(-{(|{p0,p16,p12}),((p2?p8:b1)=={p17,a5})})});
  assign y11 = ((^(~&(4'sd5)))>>>(2'd0));
  assign y12 = (-(|{{{p2,p16},(^p11)},((^p1)?{p14,p3,b2}:(p7?p4:p17)),(^{(|(^p16))})}));
  assign y13 = ((((b0!==b0)===(b2>>b0))<<({p16}<<(p16^p0)))+{2{{{1{(p0&&p13)}}}}});
  assign y14 = {((~^(((!a5)===(-4'sd2))||((-5'sd9)&(a5||a0))))>(((+a0)&&(~&b3))>={{a2,b3,p9}}))};
  assign y15 = ((|(^(p13?b4:p9)))?(~(p17?p14:p10)):$unsigned($signed((p9?p10:p13))));
  assign y16 = (((p15?a2:p2)&&(!b5))!=((-p12)?(a0!==a0):{p10,p9,b3}));
  assign y17 = $unsigned($signed((-3'sd0)));
endmodule
