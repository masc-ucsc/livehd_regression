module expression_00813(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^(~(~&(!((~&(3'sd2))||(~^(4'd3)))))));
  localparam [4:0] p1 = {2{((5'd15)&&(-4'sd2))}};
  localparam [5:0] p2 = (-2'sd0);
  localparam signed [3:0] p3 = {2{(-{1{((3'd3)^(4'd11))}})}};
  localparam signed [4:0] p4 = ((4'd0)>=(-2'sd1));
  localparam signed [5:0] p5 = (((5'sd6)!==(5'd10))/(-2'sd1));
  localparam [3:0] p6 = (5'd21);
  localparam [4:0] p7 = ((2'd2)?((-5'sd10)?(3'sd3):(-3'sd1)):{(2'sd0)});
  localparam [5:0] p8 = {{{((-3'sd2)==(3'd1))}}};
  localparam signed [3:0] p9 = (5'd30);
  localparam signed [4:0] p10 = {1{(^{2{{1{(!{1{(~|(3'd6))}})}}}})}};
  localparam signed [5:0] p11 = (((-2'sd0)%(-5'sd9))?(5'd23):((4'd10)?(4'sd5):(2'd1)));
  localparam [3:0] p12 = (~^(~|{1{(&(&{4{(~|(-2'sd1))}}))}}));
  localparam [4:0] p13 = ({4{(5'd20)}}&&(((3'sd3)>>(3'sd1))<<(5'sd0)));
  localparam [5:0] p14 = {{{(4'sd6),(2'd3),(-2'sd0)},{(5'sd11)},{(2'd2),(-2'sd0),(-5'sd1)}}};
  localparam signed [3:0] p15 = (!(|((~&((3'sd1)||(-5'sd13)))===(-((3'd5)-(4'd12))))));
  localparam signed [4:0] p16 = {(^((-4'sd5)&&(5'd18))),(^((5'd25)>>(5'sd12)))};
  localparam signed [5:0] p17 = ((5'd24)&(5'd24));

  assign y0 = (-((~|(|(~^(|(^(&(&(^(+b3)))))))))<{4{(a3+a2)}}));
  assign y1 = (5'd31);
  assign y2 = ($signed({a4})&&(-4'sd5));
  assign y3 = ((&((a3&&a1)!==(b0?a2:a4)))?({(!a1)}&(~^(p17>>b1))):((^(&b5))|(a0>>b5)));
  assign y4 = ($unsigned({{a4},(p17?a2:b4),(p12)})<<<{{(a1||p2)},(p3?b0:b5),(p12!=p8)});
  assign y5 = ((p6%p7)?(^(a4^a3)):(4'd0));
  assign y6 = (6'd2 * (p8&&p12));
  assign y7 = (|((~|p0)==(~|p9)));
  assign y8 = (~p15);
  assign y9 = {{((b5==a5)<=(b5?p11:b3))},{{(~&(p17^~p0))},(b5?p5:a4)}};
  assign y10 = {1{p5}};
  assign y11 = (((a0&&a0)|(p4||b4))&&((5'd25)<(b1>>b2)));
  assign y12 = ($unsigned((|{2{b0}}))?((a4?b4:a2)===(b1-a1)):((b4>a2)===(-a2)));
  assign y13 = (~{(($unsigned(b5)^~{p9,p12})),(+((+$signed($signed(b1))))),((~^p17)?(b4?p14:b3):(p5))});
  assign y14 = ((~&((a4==a2)===$signed((^b1))))!=={$unsigned({(b0|a4),{b2,a3}})});
  assign y15 = ({4{(p9<<<b4)}}||(-{3{(p4<b2)}}));
  assign y16 = ((a2^~p15)>$unsigned(p2));
  assign y17 = (((a3+a5)!=(4'd2 * b1))!=(6'd2 * $unsigned((a0<=b5))));
endmodule
