module expression_00170(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((6'd2 * (2'd0))?{(4'd12),(-5'sd15)}:{(4'sd7),(5'sd6),(-3'sd2)});
  localparam [4:0] p1 = ({(~^(5'd5))}>((4'd11)<(4'd3)));
  localparam [5:0] p2 = {1{(3'd4)}};
  localparam signed [3:0] p3 = (~^(!{(|({(-2'sd0),(5'sd0),(-4'sd6)}!={(4'd9)})),(+(&((!(-4'sd5))<={(2'd0),(3'd3)})))}));
  localparam signed [4:0] p4 = (2'd0);
  localparam signed [5:0] p5 = (^({((3'd0)<=(2'd0)),((-5'sd0)-(4'sd2))}<(((2'd3)!==(3'd3))&&(~(4'sd0)))));
  localparam [3:0] p6 = ((-2'sd0)<<<(3'sd2));
  localparam [4:0] p7 = ((-4'sd2)&(3'd0));
  localparam [5:0] p8 = (2'sd0);
  localparam signed [3:0] p9 = ((-2'sd1)?{1{((-4'sd3)?(5'd27):(5'd8))}}:(-2'sd1));
  localparam signed [4:0] p10 = {3{{3{(5'sd10)}}}};
  localparam signed [5:0] p11 = {3{(3'd0)}};
  localparam [3:0] p12 = (~^(~^(^(5'sd6))));
  localparam [4:0] p13 = (+{2{(-2'sd1)}});
  localparam [5:0] p14 = ((((3'd4)-(-2'sd1))?{4{(5'd26)}}:((5'd2)^~(-2'sd0)))>(4'd5));
  localparam signed [3:0] p15 = {1{{3{(4'd10)}}}};
  localparam signed [4:0] p16 = (2'd2);
  localparam signed [5:0] p17 = ((-5'sd4)?(3'd6):(5'd16));

  assign y0 = $signed((+(&(~(-p6)))));
  assign y1 = (($unsigned((~(p2?p7:a1))))?$unsigned({(&(^(p4)))}):((p0?p3:p12)?{p11}:(|a5)));
  assign y2 = (p3>>b5);
  assign y3 = $unsigned({(^($unsigned((~|(p14<<<p6)))+((b2!==b1)+(!p2)))),$unsigned({$signed({a5,p8}),{(~|(!p10))}})});
  assign y4 = (~^(&(-3'sd3)));
  assign y5 = (4'd6);
  assign y6 = (((-3'sd1)?(+((|(-3'sd1))==(|(3'd0)))):(|(3'd4))));
  assign y7 = {{(~(~^(a5==b2))),({b3,a2,b5}>=(~|a3)),{{b1,b5,b2}}}};
  assign y8 = ((5'd24)?(2'd2):{p4});
  assign y9 = {4{(p2?p8:b2)}};
  assign y10 = (((b3<b2)!==(b0>>a1))&(4'sd5));
  assign y11 = ($unsigned(p13)&(-a3));
  assign y12 = $unsigned($signed((~&(^(-(|(+(~|$unsigned(a5)))))))));
  assign y13 = (~|({(~|{a4})}));
  assign y14 = (6'd2 * (p13-p12));
  assign y15 = {{{(4'd8),{1{p4}}}},{4{p12}}};
  assign y16 = (&(~^(^(((({$unsigned((p6||b4)),(+(p16>p5))})))>=(6'd2 * (p12<=p12))))));
  assign y17 = {1{{4{(p15-p17)}}}};
endmodule
