module expression_00574(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'd3)?(4'sd0):(-5'sd12))?(5'd9):((-5'sd3)?(2'sd0):(4'sd3)));
  localparam [4:0] p1 = (((5'sd6)>=(3'd7))^~(2'd0));
  localparam [5:0] p2 = (~^(~{(+(-2'sd1)),((-3'sd1)?(4'd3):(4'd8)),(|(2'sd0))}));
  localparam signed [3:0] p3 = (+(((4'sd4)&&(2'sd0))!={(-4'sd7),(5'd26),(3'sd1)}));
  localparam signed [4:0] p4 = (4'sd7);
  localparam signed [5:0] p5 = (((2'sd0)?(4'd13):(-4'sd3))?(((5'sd0)>>(3'sd2))+(5'd6)):((2'sd0)?(5'sd15):(-2'sd1)));
  localparam [3:0] p6 = ((((3'd3)!==(3'd0))&&(|((4'sd0)<<(5'sd15))))<(|{((-3'sd0)^(5'sd15)),((2'd3)|(-2'sd0))}));
  localparam [4:0] p7 = {{2{(2'sd0)}},{2{(4'd14)}},{3{(2'd0)}}};
  localparam [5:0] p8 = {((5'd11)?(4'd2):(-4'sd1)),((-3'sd2)?(5'd12):(5'd12))};
  localparam signed [3:0] p9 = {4{((4'd1)&(2'd0))}};
  localparam signed [4:0] p10 = ((5'sd3)?(3'sd0):(-3'sd2));
  localparam signed [5:0] p11 = ((-5'sd6)!=(4'd15));
  localparam [3:0] p12 = {1{(3'd4)}};
  localparam [4:0] p13 = (((4'd2)||(4'd8))<<<((4'sd1)&(3'd0)));
  localparam [5:0] p14 = ((5'sd0)?(-4'sd2):(5'd29));
  localparam signed [3:0] p15 = {2{{1{{4{(-2'sd0)}}}}}};
  localparam signed [4:0] p16 = (&(-(2'sd1)));
  localparam signed [5:0] p17 = (((3'sd0)&(4'd4))%(2'd1));

  assign y0 = (~^(((|(~&(&b0)))===(~&(~(b4+a5))))&(!((~^(^p16))&&(p17>=b3)))));
  assign y1 = (&a3);
  assign y2 = (^(4'd1));
  assign y3 = (({4{a1}}===(b2<a2))?(4'd13):{1{(5'd15)}});
  assign y4 = (-5'sd4);
  assign y5 = ((a1&p6)<<(b3^p17));
  assign y6 = (~&(({b3,p9})?(~(~|{b5,p17,b0})):($signed(p1)!=(~a5))));
  assign y7 = (((^{(p11^~a1),{2{a1}}})^(5'd2 * (!(a1<<p14))))<={(~|(|{1{{a5}}})),{(p13&b3),(~|b3),{p0}}});
  assign y8 = ({2{((b3===b0)||(5'd2 * p14))}}==((b4>=b3)?({a4,b2}):(-(-5'sd6))));
  assign y9 = (p11^a2);
  assign y10 = (!(6'd2 * (p12|p7)));
  assign y11 = {4{{1{b4}}}};
  assign y12 = (6'd2 * (p8/p1));
  assign y13 = (&(&{(!(~^{p8,p5})),{(~&b2),{b4,a5},(~|b5)},(|{(!b1),{b0}})}));
  assign y14 = (6'd2 * {b1,p13,a1});
  assign y15 = (((a3!==b5)?(p6<<a1):(b4|p9))?((p2/b2)<<<(a1?p11:p6)):((a1^b1)!==(a3&&b5)));
  assign y16 = (&((|(|((-2'sd1)?({(a0>>b5)}!={b1,p6}):(2'sd0))))));
  assign y17 = (((-5'sd0)+(-4'sd6))>=((p3?p13:p9)?(4'd10):(3'sd2)));
endmodule
