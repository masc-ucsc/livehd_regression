module expression_00772(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'd3)^~(-5'sd10))/(4'd9))>>(((2'd1)==(5'd4))+((3'd1)<<(5'd13))));
  localparam [4:0] p1 = (^(~&(~(-(^(|(3'sd3)))))));
  localparam [5:0] p2 = {4{{4{(3'sd2)}}}};
  localparam signed [3:0] p3 = ((2'd2)||(-4'sd7));
  localparam signed [4:0] p4 = (+(~(~|(~^(&(~(~|(2'd2))))))));
  localparam signed [5:0] p5 = ((((4'd0)^(5'd26))^~(2'd2))<((~^(5'd19))<(!(|(4'sd0)))));
  localparam [3:0] p6 = {(((-3'sd3)>>(-3'sd3))<((4'sd3)?(-4'sd3):(5'd0)))};
  localparam [4:0] p7 = (!{1{(-{{{4{(5'd22)}}},((~^(-4'sd6))==((-5'sd0)||(4'd13)))})}});
  localparam [5:0] p8 = {4{(4'd4)}};
  localparam signed [3:0] p9 = (4'd14);
  localparam signed [4:0] p10 = (-5'sd3);
  localparam signed [5:0] p11 = (-3'sd1);
  localparam [3:0] p12 = (((3'd4)==(-5'sd3))-(2'sd1));
  localparam [4:0] p13 = {((-5'sd12)<(3'd5)),(~(-2'sd1))};
  localparam [5:0] p14 = (((~(-2'sd0))?(^(4'd11)):((2'd2)<<(-3'sd0)))<<<{((4'd10)<<(3'd0)),(~(|(3'd0)))});
  localparam signed [3:0] p15 = (|(~&(&(+(!({4{(5'd10)}}^~(-({1{(3'd7)}}==((3'sd3)===(3'd3))))))))));
  localparam signed [4:0] p16 = (^(((5'd18)||(2'sd0))^((-4'sd5)>>(-2'sd1))));
  localparam signed [5:0] p17 = (((4'd9)?(5'd24):(5'sd4))?(6'd2 * ((2'd1)&&(4'd11))):((5'd20)?(-3'sd2):(2'd0)));

  assign y0 = (4'sd5);
  assign y1 = ({p0}+{1{p3}});
  assign y2 = {{p7,p4,a1},((p12?p15:p2)-(^a3)),{{p14,p8}}};
  assign y3 = $unsigned((p16>=p3));
  assign y4 = (a2===a5);
  assign y5 = (~|{(~&{4{p8}}),{(~^a0),{b1,p4},{1{b3}}},(~|{(p17+b3)})});
  assign y6 = (((-3'sd0)-(~|p11))<<(!((a4<b5)-(~^p12))));
  assign y7 = (4'sd1);
  assign y8 = (~|((~(!(p16-p8)))&&(2'sd0)));
  assign y9 = (((p7^p10)|(p5|p14))?((p14<<<p7)<<<(b3^p15)):((p6<<p0)>>>(p17>=p3)));
  assign y10 = ((+{((^((|(!($signed(a5)-$unsigned(a2))))==(~&({p10,a3,a2}>=$unsigned((&b3)))))))}));
  assign y11 = ({2{(2'sd0)}}^~{2{{{b2,p2},{2{p4}}}}});
  assign y12 = {3{(-((b1|p16)||(a3<b1)))}};
  assign y13 = ((b5<a1)!=(b5===b0));
  assign y14 = (4'd5);
  assign y15 = ((((4'd1)&&$unsigned({b4,b3,b5})))<({a5,p11,p2}>(2'sd1)));
  assign y16 = $signed((3'd6));
  assign y17 = {2{({b5,b0}-(p16>=a5))}};
endmodule
