module expression_00921(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'sd7)?(-2'sd1):(2'd2));
  localparam [4:0] p1 = (^{((^(|(2'd2)))?((5'sd10)|(4'sd2)):(^(~|(-2'sd1))))});
  localparam [5:0] p2 = {{4{(5'd10)}},{(-2'sd1),(5'd22),(3'sd0)},{1{(5'sd0)}}};
  localparam signed [3:0] p3 = (&(-{(~^(~|{3{{3{(4'd13)}}}}))}));
  localparam signed [4:0] p4 = (!{2{((~&(-4'sd1))?(3'sd0):(~&(2'sd0)))}});
  localparam signed [5:0] p5 = {{(3'd1),(2'd1),(5'd2)},((4'd15)&&(2'sd1)),((-5'sd0)>=(4'd12))};
  localparam [3:0] p6 = (|(3'sd3));
  localparam [4:0] p7 = (3'd0);
  localparam [5:0] p8 = (-(5'd18));
  localparam signed [3:0] p9 = (&((-(((5'd11)<<(-5'sd10))>=((4'sd6)>>(-4'sd0))))&(((2'd0)<<<(3'sd2))!==(~^(4'sd4)))));
  localparam signed [4:0] p10 = ((2'd1)?(4'd11):(2'd1));
  localparam signed [5:0] p11 = ((-3'sd2)==(4'sd0));
  localparam [3:0] p12 = {{{(5'sd2),(4'd13)},{(2'd1),(4'd2),(2'd3)},((2'd3)-(-5'sd3))},{(5'd2 * ((3'd4)-(2'd3)))}};
  localparam [4:0] p13 = {2{(2'd0)}};
  localparam [5:0] p14 = (((4'sd6)<(5'd21))?(6'd2 * (5'd30)):((-4'sd0)<<(5'd17)));
  localparam signed [3:0] p15 = {(-2'sd0),(2'd1)};
  localparam signed [4:0] p16 = ((-5'sd8)&&(4'd2));
  localparam signed [5:0] p17 = (~&(~&({(2'sd0),(-2'sd1),(-2'sd0)}>>>(+(5'd0)))));

  assign y0 = $unsigned(($unsigned((p5||p14))||$signed($signed((p11||a1)))));
  assign y1 = (!{{p2}});
  assign y2 = ($signed(((b2>>>b5)?{a2,a1}:(a0)))?({a3,b0}>>>(p5?a2:b3)):{(a3<<a2),(a3>=b0)});
  assign y3 = ((4'd15)/p3);
  assign y4 = {1{{2{(^((p15?p4:p15)?(^p13):(!p11)))}}}};
  assign y5 = (($unsigned((a1?a2:p15))<=(b1/b5))?((b1>b0)!==(b3||b5)):(!(~^((a3+p14)<<$signed(p5)))));
  assign y6 = ($signed((((!a0)^~(b1))&(2'd1)))!==((4'sd2)));
  assign y7 = ({2{(5'sd14)}}?{2{{1{(b3?a5:b1)}}}}:{({3{b2}}?(2'd3):(-3'sd1))});
  assign y8 = (((-3'sd1)^{1{b5}})>>>(^(~|(b5||a0))));
  assign y9 = (~^(&(~((p16?p9:p11)?(~|a5):(a0>b0)))));
  assign y10 = (+((a1?p8:a5)%p5));
  assign y11 = (2'd1);
  assign y12 = ((((a0+a5)^(a5===a4))!==((a4>>>b3)>>>(b3?b3:a3)))<=(2'd3));
  assign y13 = $unsigned($unsigned(((((((a3<<<p16)|$unsigned(p9))<<(^(a1-a2))))))));
  assign y14 = (|(|(|(-(|(~|(|a4)))))));
  assign y15 = (-$signed(((~|(~^(^(-4'sd0))))<<(-5'sd12))));
  assign y16 = (+(~|(((b3-a0)?(b3?b1:a4):(a1==a2))?((a2+b0)?(&b3):(^p2)):(-(a4?a2:a2)))));
  assign y17 = ($unsigned((-$unsigned(b3))));
endmodule
