module expression_00111(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{(-4'sd3)}}||{(4'sd6),(-4'sd7)});
  localparam [4:0] p1 = (((3'd5)^(4'd9))*((3'd1)||(-3'sd0)));
  localparam [5:0] p2 = (((5'd22)?(-4'sd7):(3'sd3))?((3'sd1)?(-2'sd0):(-5'sd4)):((5'd29)?(3'sd2):(3'd1)));
  localparam signed [3:0] p3 = (~|((!(~&(&(-3'sd1))))+((+(5'd13))==((4'd1)<(3'sd2)))));
  localparam signed [4:0] p4 = (-3'sd2);
  localparam signed [5:0] p5 = (6'd2 * ((5'd15)>>(4'd13)));
  localparam [3:0] p6 = {1{(4'd1)}};
  localparam [4:0] p7 = (((2'd0)?(-2'sd0):(5'sd3))?((2'd1)>>(4'sd2)):((5'sd12)?(3'sd3):(5'sd3)));
  localparam [5:0] p8 = (((-5'sd10)>>(2'd1))^~((-3'sd2)<(5'd31)));
  localparam signed [3:0] p9 = ((2'd2)===(|(((-3'sd1)==(3'd1))+(2'd1))));
  localparam signed [4:0] p10 = (4'sd5);
  localparam signed [5:0] p11 = (((2'd0)?(-4'sd1):(2'd3))?((-4'sd6)||(4'sd3)):((2'sd1)?(5'sd6):(-5'sd9)));
  localparam [3:0] p12 = (((3'sd3)<=(2'd0))+{4{(5'd18)}});
  localparam [4:0] p13 = {{(3'sd1),{1{{(5'd30),(-2'sd1),(5'd17)}}}}};
  localparam [5:0] p14 = (({3{(4'sd5)}}?{1{(4'sd6)}}:((5'd21)-(3'd2)))|(|{3{((2'd3)>>(5'd21))}}));
  localparam signed [3:0] p15 = ((2'd3)>(5'sd6));
  localparam signed [4:0] p16 = (2'sd0);
  localparam signed [5:0] p17 = (~^(~|(4'd9)));

  assign y0 = {p12,b2,p10};
  assign y1 = ((p6<<p14)?(p10>=p12):(b2<a1));
  assign y2 = ((-4'sd6)<=((-4'sd4)?(4'd1):(-5'sd1)));
  assign y3 = (~^((a3===b4)*(p2-p10)));
  assign y4 = {1{((($unsigned(a4)!==(a2))==((p10>=b5)^~(b4^p10)))<<(+((5'd2 * b0)||((p16&&p12)))))}};
  assign y5 = (&(!{(~|(p5?p11:p12)),(p6?p4:p11),(~|(p7?p15:p13))}));
  assign y6 = ((p6|p0)|(p7&p4));
  assign y7 = ((6'd2 * (!{1{b0}}))|(^{2{(!(&b0))}}));
  assign y8 = $unsigned((p14?p5:p17));
  assign y9 = (-(~(^{$unsigned({(5'd8),(|a1)}),(^$unsigned({(5'd21),(2'sd0)})),{{p3,p5},$unsigned($unsigned(b1))}})));
  assign y10 = (p2^~p1);
  assign y11 = {(a1===b1),{p16,p14,p16}};
  assign y12 = ({4{a1}}?((!p13)||(p2!=a2)):(^(b3?p2:p5)));
  assign y13 = {1{(a3^~a1)}};
  assign y14 = ({1{((p11?p16:p1)?(p5?p13:b5):{4{p14}})}}>>>(((b3?b0:p15)&(a0!=p9))|((p13!=p11)?(p17>p8):(p8+p17))));
  assign y15 = $unsigned((~&($signed((-((p6>>>p10)))))));
  assign y16 = (5'd2 * (a0?b1:p7));
  assign y17 = (((p1||a1)^(p5?b3:b2))?(^{{b1,b1,p13}}):((!p11)?{b1,p2,p0}:(b0?p6:a1)));
endmodule
