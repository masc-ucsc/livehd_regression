module expression_00976(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (6'd2 * ((4'd1)-(4'd5)));
  localparam [4:0] p1 = ((-2'sd0)?{((-4'sd0)?(-4'sd4):(3'd2))}:{{(&(5'd5))}});
  localparam [5:0] p2 = {1{(^((-{4{(3'd3)}})^{1{(^((3'd1)^~(-2'sd1)))}}))}};
  localparam signed [3:0] p3 = {(2'sd1),(-2'sd0)};
  localparam signed [4:0] p4 = (~&((&(((4'd8)===(5'd16))%(3'd7)))==(^(|(~&((-3'sd1)<=(2'd1)))))));
  localparam signed [5:0] p5 = (((2'd1)>=(-5'sd0))>={2{(2'd2)}});
  localparam [3:0] p6 = ((-4'sd0)?(3'd3):(-2'sd0));
  localparam [4:0] p7 = (((^(-4'sd2))?{(2'd0),(2'd0),(-5'sd7)}:{(3'd1),(2'd0)})!==(5'd19));
  localparam [5:0] p8 = (2'sd1);
  localparam signed [3:0] p9 = ((+(&(!(~|(4'sd2)))))!=(~&(!((3'd3)?(-4'sd1):(5'd1)))));
  localparam signed [4:0] p10 = {2{{(5'd4),(-5'sd15)}}};
  localparam signed [5:0] p11 = {((((4'sd2)&(-2'sd0))&((5'd15)^~(-5'sd1)))===(((5'd5)!=(3'sd3))|((-3'sd2)&&(5'd8))))};
  localparam [3:0] p12 = (((5'd22)<(2'd0))<{3{(5'd18)}});
  localparam [4:0] p13 = (((|(-(-5'sd10)))&((5'sd0)>(-4'sd2)))<<(((-2'sd0)||(3'sd3))<((5'd27)^(5'd21))));
  localparam [5:0] p14 = (~^({2{{4{(3'd2)}}}}>=(|{1{(~|{3{(5'd10)}})}})));
  localparam signed [3:0] p15 = (^(5'd8));
  localparam signed [4:0] p16 = {(((|(2'd0))?(^(-4'sd6)):((5'sd5)+(4'd8)))?(&{((4'd2)?(3'd0):(2'd0)),((3'd3)===(3'd7))}):({(3'sd1),(-2'sd1)}?((4'd7)<(-4'sd6)):((2'sd1)?(2'd0):(-4'sd1))))};
  localparam signed [5:0] p17 = (5'd28);

  assign y0 = {1{({b1,a1,p4}^~(b2?p2:p17))}};
  assign y1 = {{((^(&b3))<<(b0>>>p14)),((p1!=p2)<(&(~^a0))),(&({a4}-{b2}))}};
  assign y2 = {3{$signed((&p6))}};
  assign y3 = (&(~(&(^((2'd2)+(-5'sd13))))));
  assign y4 = (((~&p14)?{b4,p13,b2}:(3'sd3))?((^a3)?(-4'sd5):{p10,a1,a5}):(-4'sd7));
  assign y5 = $unsigned((((-2'sd1)-((~^a4)>=(a0-a2)))==(((p13&&a1)<<<(p1<<a5))>=(5'd1))));
  assign y6 = {(p13&&p13),{p12,p15}};
  assign y7 = (-(~^(~&((-3'sd0)>=(((p15!=p7)&(a0==p6)))))));
  assign y8 = $signed({1{$unsigned((-5'sd3))}});
  assign y9 = ((~^{(~p9),{a3,a0},{a5}})<<<{(b1>=a4),(b4>>b5),(a3-a1)});
  assign y10 = (({1{{3{a5}}}}||((a1>>>p5)==(p0&a5)))<<<((^((a2>a3)))!==($unsigned(b5)!=={3{b1}})));
  assign y11 = ((|((+p7)|(p15%p16)))!=((a4<<<p5)>(p12/p14)));
  assign y12 = ((!(~^((p10?a2:b2)?(a2>>>b4):(~|p17)))));
  assign y13 = {{p7,p11},$signed(p11),(a2<<<a1)};
  assign y14 = (5'd2 * (4'd2));
  assign y15 = ((-3'sd3)<<<({p2,b0,b4}>>>((~&a3)>>>(a5&&b2))));
  assign y16 = (~{4{p14}});
  assign y17 = ((4'd2 * p1)?(+(-p16)):$unsigned((p6/p15)));
endmodule
