module expression_00506(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(~|((-4'sd2)!==(-3'sd0)))}};
  localparam [4:0] p1 = (+{4{(-4'sd4)}});
  localparam [5:0] p2 = (+(3'd5));
  localparam signed [3:0] p3 = {1{(|((~|(4'd13))+((2'd1)<<<(4'sd2))))}};
  localparam signed [4:0] p4 = (~^(~&{2{{3{((3'd5)===(4'd15))}}}}));
  localparam signed [5:0] p5 = (~&(((^(-4'sd5))||(|(4'sd1)))^(!(~^((2'd2)+(4'sd5))))));
  localparam [3:0] p6 = {1{((((3'd5)^(4'd5))>>>(~|(3'd3)))!=((-(~|(-3'sd3)))==={2{(2'd3)}}))}};
  localparam [4:0] p7 = (|((((-3'sd3)>>(2'd0))=={(-2'sd0),(3'd3)})>>>(+{(3'sd2),(4'd2),(-4'sd7)})));
  localparam [5:0] p8 = (~|{(!(|{(-3'sd1)})),(~&(!{(3'sd3),(4'd2),(-4'sd7)})),(2'sd1)});
  localparam signed [3:0] p9 = {4{{2{(2'sd1)}}}};
  localparam signed [4:0] p10 = (~(|(~&{{({(4'd13)}|{4{(3'd0)}}),(((2'd3)?(3'sd0):(3'd7))<=(&(4'd2)))}})));
  localparam signed [5:0] p11 = (~&((^(-4'sd4))<(-(4'sd0))));
  localparam [3:0] p12 = {2{(4'd14)}};
  localparam [4:0] p13 = (|((2'sd0)!==(-3'sd1)));
  localparam [5:0] p14 = ((~^(4'd13))>>>(~&((&(3'd1))?(~|(4'sd7)):(!(-3'sd0)))));
  localparam signed [3:0] p15 = ((((3'd1)!==(3'd4))>>((-4'sd6)?(2'd3):(-3'sd1)))|(((-2'sd0)?(5'd27):(3'd2))<<((5'd0)==(5'd24))));
  localparam signed [4:0] p16 = (~|(~&((((3'd0)-(3'd6))===((4'sd1)?(2'sd1):(-2'sd1)))?(((5'd0)<(3'd2))/(-2'sd1)):((-5'sd0)?(3'd0):(3'd6)))));
  localparam signed [5:0] p17 = {(((4'd10)>=(2'd1))^((4'sd6)^(-3'sd1))),(((5'sd11)>>(-2'sd1))<=((-2'sd0)<<(4'd13))),((3'd4)?(5'd30):(4'sd3))};

  assign y0 = (~|(~|((a2?b3:a3)==(+b5))));
  assign y1 = ({4{$unsigned(a5)}});
  assign y2 = (((2'sd1)>>(4'd15))?{2{(2'sd1)}}:{4{p6}});
  assign y3 = {(a2<b0),(5'd2 * a0)};
  assign y4 = {((p9?p4:p17)?{p5,p4}:(2'd2)),(2'd1),(4'd2)};
  assign y5 = (((b3!=b4)!={b1,b2})<<<$unsigned({(b5|p7),{2{p13}},$signed(b5)}));
  assign y6 = (~(~(-(4'd4))));
  assign y7 = (^((~(~|(-4'sd5)))<=(&((p2!=p13)<<(5'd7)))));
  assign y8 = (4'sd1);
  assign y9 = (-((&(|(p14<<<b3)))<=((~|p11)/b2)));
  assign y10 = {1{((4'd5))}};
  assign y11 = {{{b2,b5},{a2,a0,b2},(b2!=b3)},{{(4'd2 * {(a1!==a1)})}}};
  assign y12 = (((~&(~((|(~((3'd4)))))))));
  assign y13 = (~&(~(!{4{(&{a3})}})));
  assign y14 = (^(+(+(~&(|{b1})))));
  assign y15 = (~&{3{(-(2'sd0))}});
  assign y16 = {{(p15?p1:p16)},((^p0)?(~p7):(~&p10)),{(p6?p13:p13),(p14?p12:p7),(!p11)}};
  assign y17 = (3'd3);
endmodule
