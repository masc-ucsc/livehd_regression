module expression_00503(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {({(5'sd14)}^((-3'sd2)<=(5'd17))),(~{{1{{3{(5'sd2)}}}}}),({(5'sd5),(-4'sd5),(2'd3)}<{1{(5'sd5)}})};
  localparam [4:0] p1 = ((6'd2 * ((4'd8)>>>(3'd4)))<<<(&({(-4'sd5),(3'sd1)}^~((-4'sd4)>=(2'd3)))));
  localparam [5:0] p2 = {(~^(3'd6)),(5'd28),(-(3'd3))};
  localparam signed [3:0] p3 = (^(+((5'd27)?(2'sd0):(4'sd7))));
  localparam signed [4:0] p4 = ({3{(5'd11)}}?(!(4'sd3)):((5'd15)?(3'd4):(5'sd10)));
  localparam signed [5:0] p5 = {(2'd2),(2'sd1),(2'sd0)};
  localparam [3:0] p6 = (&(2'sd1));
  localparam [4:0] p7 = ({2{(2'd3)}}?((-3'sd0)?(2'sd1):(3'd2)):((2'd1)>=(5'sd1)));
  localparam [5:0] p8 = (3'd0);
  localparam signed [3:0] p9 = (|(4'd9));
  localparam signed [4:0] p10 = ((|(-(2'd2)))!=((4'sd3)*(2'd3)));
  localparam signed [5:0] p11 = (-(-(+(~&{3{(((4'd6)!==(-3'sd1))=={4{(-3'sd1)}})}}))));
  localparam [3:0] p12 = (~(~^(2'd3)));
  localparam [4:0] p13 = (3'd6);
  localparam [5:0] p14 = (((-4'sd1)?(3'd5):(-4'sd3))&((4'd7)^~(4'd15)));
  localparam signed [3:0] p15 = (!{2{(+{{1{(4'd12)}},(~(5'sd5)),((-3'sd1)?(5'sd12):(5'd18))})}});
  localparam signed [4:0] p16 = (((-4'sd6)>=(-2'sd0))<=((3'sd2)&(2'd0)));
  localparam signed [5:0] p17 = {1{{(~|((3'sd3)<<(5'd15))),{(-2'sd0),(-3'sd2),(-2'sd1)}}}};

  assign y0 = {(~{4{{3{p11}}}}),(&{(b2^~p16),{p16,p2,p3}})};
  assign y1 = (({3{b3}}&&({2{a3}}))?(((4'd5))<<(a2?p2:b5)):(-3'sd0));
  assign y2 = $signed((((a0<<<b0)?(b0<<<a5):(a0<=a3))<((~^a1)?(b5==a0):(5'd26))));
  assign y3 = ((-(((a2&&a1)==(~|a1))===(&(&(a2!=a1)))))||(((~|b2)+(|p10))==(p12?p12:b3)));
  assign y4 = ($signed($unsigned(((~&$signed((b3===b4)))<<((~&a0)||$signed(a5)))))<<<$signed((($unsigned(a0)<<<(b1||b4))<{$unsigned($unsigned(b4))})));
  assign y5 = ((+{1{(b2|b0)}})&(!(2'd0)));
  assign y6 = {(|(|((~(~^{(!a5),(&p6)}))?(&{(+(p0?p17:p8))}):((p4?p4:p9)?(!p9):(+p7)))))};
  assign y7 = (p15?p9:p17);
  assign y8 = ($signed({2{{p9,b3}}}));
  assign y9 = ((6'd2 * b0)?(b5||b0):(~p9));
  assign y10 = ({b0}<(b1&&a5));
  assign y11 = (~{{{(~(+{b2,b4,a3})),(~&{b3,b1})},{(&{{(^b3),(~b5),{a1,b4}}})}}});
  assign y12 = (b1&&p17);
  assign y13 = {(|a1),(a1)};
  assign y14 = (((b1!==a0)<<<(3'd2))?(2'd0):((p8?p4:p16)?(-2'sd1):(p8?p12:p5)));
  assign y15 = (^({(+p12),(^p15)}<<((~|a0)>(a2||a4))));
  assign y16 = ((-{a5,p7})!=(4'd10));
  assign y17 = (!(!(+(5'd7))));
endmodule
