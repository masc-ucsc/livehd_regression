module expression_00238(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd0);
  localparam [4:0] p1 = {(((3'd7)&(4'd0))>>(3'd5)),((2'd3)||(2'd0))};
  localparam [5:0] p2 = {2{(6'd2 * (~(&(2'd2))))}};
  localparam signed [3:0] p3 = {{(-(4'sd2)),{(2'd3)},(|(4'sd5))},(&(+{(~|{(2'd3),(2'sd1),(-2'sd0)})}))};
  localparam signed [4:0] p4 = {2{{(3'd3)}}};
  localparam signed [5:0] p5 = (4'd10);
  localparam [3:0] p6 = (4'd2 * (-((5'd17)?(3'd1):(4'd6))));
  localparam [4:0] p7 = (-4'sd4);
  localparam [5:0] p8 = (4'd15);
  localparam signed [3:0] p9 = ((~(5'd30))<<<(((4'sd5)-(5'sd9))==={(4'd13),(4'd0),(4'd8)}));
  localparam signed [4:0] p10 = (((3'd1)||(2'd3))/(5'd1));
  localparam signed [5:0] p11 = (((4'd5)===(3'd4))||((3'd5)<<<(5'd20)));
  localparam [3:0] p12 = (2'd1);
  localparam [4:0] p13 = {1{((2'sd0)^~(((-4'sd5)>>(3'd0))==(-3'sd2)))}};
  localparam [5:0] p14 = ((-(!({(-4'sd2)}<(~&(4'd6)))))>=(4'd2 * (~|((5'd10)>=(5'd2)))));
  localparam signed [3:0] p15 = ((((2'd0)?(2'd1):(4'd13))*((5'sd0)<<(-3'sd0)))?(((3'sd0)^(4'd4))^~((-2'sd1)-(2'sd1))):((5'd2 * (2'd2))^~((-4'sd2)^(-5'sd12))));
  localparam signed [4:0] p16 = ((2'd1)?(5'd5):(3'd6));
  localparam signed [5:0] p17 = (-4'sd4);

  assign y0 = $signed({$signed({3{{p5}}}),({1{(p13-p7)}}>={1{$signed(p2)}})});
  assign y1 = ((3'd5)==(&(!((~|(p11>a3))>=((p15&&p6)^~(-2'sd0))))));
  assign y2 = (4'd2 * (!a1));
  assign y3 = (((-(-(+p15)))^~(p7?p13:a2)));
  assign y4 = ((6'd2 * (b1<=a0))!==((5'd2 * (3'd2))<((3'd6)&(b3!==a1))));
  assign y5 = (p7?p6:p15);
  assign y6 = $signed(p16);
  assign y7 = (((p6?a0:b5)==(~&p12))?((a5&&p3)?(~^p13):(a0?b1:p12)):((a5?a1:b0)?(b0>=b5):(p10?p9:b0)));
  assign y8 = (({1{{2{a4}}}}>(a2^b4))!=={3{{4{b2}}}});
  assign y9 = {4{(b3+b3)}};
  assign y10 = $signed((((p13>=b3))<<<((a1?a4:b2)^{2{a1}})));
  assign y11 = (~&a2);
  assign y12 = (~((-(p12+p13))&&((p9>=b1)&&(4'd1))));
  assign y13 = (((~^b5)?(5'd1):(b5==b4))?(~(-3'sd1)):(^{3{(b4?a3:b0)}}));
  assign y14 = (^((b0/b3)/a2));
  assign y15 = (a4<a2);
  assign y16 = ((3'd1)?(p14&a1):(a5^~p13));
  assign y17 = ((a0?a5:a1)?$unsigned((b3?p6:a2)):(b2?a0:b2));
endmodule
