module expression_00831(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{(3'sd1)}}<={4{(4'd12)}});
  localparam [4:0] p1 = ((~(5'd2 * ((2'd3)>>>(2'd0))))>=(~|(~(+(((3'd6)^(-2'sd1))!=(-(4'sd3)))))));
  localparam [5:0] p2 = (&(^(((3'd5)>>>(-3'sd2))<<((2'd0)+(2'd0)))));
  localparam signed [3:0] p3 = (2'sd1);
  localparam signed [4:0] p4 = (((2'd2)<<<(|((2'd1)^(5'd22))))>=(((4'd2)||(-4'sd4))?((2'd1)%(2'sd0)):((4'd4)<<(-5'sd4))));
  localparam signed [5:0] p5 = ((~&{((4'd13)-((3'd0)-(-4'sd2)))})&((3'd5)!={(3'd4),(-5'sd10),(5'sd4)}));
  localparam [3:0] p6 = (-((|{((2'sd0)?(5'd25):(5'd25))})?(((5'd30)-(5'd2))&&(~&(5'sd10))):(&{3{(3'sd2)}})));
  localparam [4:0] p7 = {((~(5'd14))?((4'd9)<(4'd11)):((2'd0)!=(3'd1))),(2'd2),(~&((3'd1)?(4'sd7):(-5'sd6)))};
  localparam [5:0] p8 = {(^(~(5'sd11))),(((3'd2)?(3'd1):(3'sd2))>(2'sd0))};
  localparam signed [3:0] p9 = ((((4'd15)||(2'd3))^~((2'd2)>(5'sd4)))===(!((2'sd0)?(-2'sd1):(4'd0))));
  localparam signed [4:0] p10 = (~^((5'd26)<<(5'd6)));
  localparam signed [5:0] p11 = (|(({3{(4'd11)}}<<<(2'sd0))==({2{(4'd7)}}^(2'sd0))));
  localparam [3:0] p12 = ({2{(3'sd3)}}?((2'd1)?(-5'sd7):(4'd9)):(&(^(5'd2))));
  localparam [4:0] p13 = (3'sd0);
  localparam [5:0] p14 = ((4'd2 * (5'd26))<<<(!{4{(-4'sd0)}}));
  localparam signed [3:0] p15 = ((4'd15)^~{2{(5'sd12)}});
  localparam signed [4:0] p16 = ((5'd2 * (3'd2))<=((4'd3)+(2'd2)));
  localparam signed [5:0] p17 = (&(-4'sd2));

  assign y0 = ((p3>p0)*(a3!==b0));
  assign y1 = (+((+((6'd2 * b2)===(b4&b2)))>>{(-b1),{a3,a3},(!b3)}));
  assign y2 = (($unsigned(b2)-(p6<=p15))?(5'sd2):(2'sd0));
  assign y3 = {(-2'sd1),{(p3>>a4),(4'sd0),{a0}},(-{4{(5'd2 * a2)}})};
  assign y4 = (b1!==a0);
  assign y5 = ((~&$signed((~$signed($signed(b4)))))>=((~{(~&p7),(~|a1)})));
  assign y6 = (p9>=p2);
  assign y7 = ($unsigned(((((-3'sd1))|(-5'sd5)))));
  assign y8 = ((~&(-((6'd2 * p13)+(a5>=p4))))<<(-(~(-(p7==b5)))));
  assign y9 = ((|{2{(5'd25)}})^(~^($signed((2'd1))>(3'd4))));
  assign y10 = (~|(!{(((b5>p11)^~(-3'sd0))&(3'd7)),{(6'd2 * a1),{a3,b2},$unsigned((p12|b4))}}));
  assign y11 = ((-{1{(b4<<p9)}})||$unsigned({1{(a2|p11)}}));
  assign y12 = (&((~&(b1?p17:b3))?((~^a2)!==$unsigned(a2)):(~{{b1},{a1,p5}})));
  assign y13 = {(p17||p13)};
  assign y14 = {4{(a1^~a0)}};
  assign y15 = ((((p0<<<a3)!=(&b1))+{(~^p1),(p1>p7)})+(((~|p10)&(p14&&p15))!={{(p17<p6)}}));
  assign y16 = (((b4!=b0)||(+(a4?b0:a4)))?((+(a1^~b5))^(|{b1,b5,a0})):((-{b0,a0})&(a3&&a1)));
  assign y17 = {({(5'd24)}^(b0>p17)),(2'd1),{(p10&p0),(p5>p4)}};
endmodule
