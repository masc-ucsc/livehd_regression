module expression_00674(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(3'sd1),(3'd5)},(~((3'd0)!=(2'd1)))};
  localparam [4:0] p1 = {2{(|(~|{3{((-4'sd4)^(-4'sd7))}}))}};
  localparam [5:0] p2 = ((~^((4'd0)!=(4'd4)))+{(5'd31),(4'd14),(-4'sd4)});
  localparam signed [3:0] p3 = {{(5'd28),(5'sd14),(-2'sd0)}};
  localparam signed [4:0] p4 = ((((3'd1)%(-2'sd0))||(3'd3))>>>(4'sd6));
  localparam signed [5:0] p5 = ({4{(-2'sd0)}}?((-2'sd1)?(-5'sd15):(-2'sd0)):((4'sd1)?(5'd7):(4'd5)));
  localparam [3:0] p6 = (|(~|(&{{(4'd13),(5'sd2)},{(-4'sd2)},(!(3'd4))})));
  localparam [4:0] p7 = {((-3'sd1)||(~|((2'd2)?(4'sd6):(5'd10))))};
  localparam [5:0] p8 = (~&(-4'sd6));
  localparam signed [3:0] p9 = {3{(5'sd1)}};
  localparam signed [4:0] p10 = {1{(-3'sd1)}};
  localparam signed [5:0] p11 = (-5'sd11);
  localparam [3:0] p12 = ((-3'sd1)&(5'sd14));
  localparam [4:0] p13 = {(({(-2'sd0)}>>(-(3'sd1)))?({(4'd12),(-4'sd5),(4'sd0)}^(+(3'd6))):(~&{(3'sd1),(3'sd0),(3'sd2)}))};
  localparam [5:0] p14 = ({(3'sd1)}>={2{(-4'sd2)}});
  localparam signed [3:0] p15 = {2{{1{{(-4'sd7),(2'd0),(3'sd3)}}}}};
  localparam signed [4:0] p16 = {{(-((2'sd1)!==(4'd1)))}};
  localparam signed [5:0] p17 = (5'd5);

  assign y0 = (((p11>>p9)%a2)<=((a5-p12)<=(p7/a0)));
  assign y1 = $unsigned({(4'd2),(b0<b0)});
  assign y2 = (~&((|(~({a0}<<<{a1})))<=({p7,b1}?{a3,b0,a2}:(|p7))));
  assign y3 = (($signed((p12/p10)))>(|($signed((p16!=p1)))));
  assign y4 = (p4<<b5);
  assign y5 = {a2};
  assign y6 = (~(-(~((((a4>b1)===(a5))|(!(&(p14-p17))))))));
  assign y7 = ((~&($unsigned((~&(-$signed((b5?b5:b4)))))))===((b4?b1:b1)<=$signed((b1^~b2))));
  assign y8 = {{({2{p0}}^~(p16<=p1))},{{3{p7}},(2'd0)}};
  assign y9 = {2{{(b0!==a3),(p12<<p14),(p11&p4)}}};
  assign y10 = {2{{1{(^p2)}}}};
  assign y11 = (((p17>=p11)-(a3?p17:p17))<<((b2&&p13)?(b5?p12:p15):(p14^~p1)));
  assign y12 = (((b2>>>b4)?(&(a1<<<b5)):(!(b0!==a2)))||({(-3'sd2)}?(p17?a4:b1):(4'd12)));
  assign y13 = (&(6'd2 * (|$unsigned(p13))));
  assign y14 = ((~&(a0?b0:b0))^~$unsigned($signed((!(p7>>b2)))));
  assign y15 = (+({p1,p6,p12}?{(p11<<a1)}:((~|a5)!==(b1))));
  assign y16 = {3{$unsigned(b3)}};
  assign y17 = (6'd2 * (~&$unsigned(a2)));
endmodule
