module expression_00518(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{(~&{4{(4'd1)}})}}};
  localparam [4:0] p1 = (^(~&(^(!(4'sd0)))));
  localparam [5:0] p2 = ((5'd5)==(-2'sd0));
  localparam signed [3:0] p3 = {{1{(2'sd0)}}};
  localparam signed [4:0] p4 = (+(3'd5));
  localparam signed [5:0] p5 = ((((4'sd3)^~(-3'sd2))+(~(6'd2 * (3'd4))))<=(((4'd8)==(2'd3))<<<((3'd4)==(3'd7))));
  localparam [3:0] p6 = (|{(!(~&(~((5'd7)?(3'sd0):(-2'sd1)))))});
  localparam [4:0] p7 = (({(-2'sd0)}>>>{(-5'sd10),(2'd0)})+((!(3'd5))|((2'd1)==(-3'sd1))));
  localparam [5:0] p8 = ((((3'd4)?(3'd5):(-4'sd6))===((3'd2)&&(3'd5)))<(((4'd13)|(4'd12))*((2'd2)>(3'd6))));
  localparam signed [3:0] p9 = (((5'sd4)?(5'sd1):(3'sd1))?((+(3'd6))-(|(3'sd0))):((5'd13)&&((2'd2)>>(5'sd8))));
  localparam signed [4:0] p10 = ((-2'sd1)!={3{(~|(-5'sd1))}});
  localparam signed [5:0] p11 = (4'd2 * {2{(2'd3)}});
  localparam [3:0] p12 = ((((5'd23)%(2'd3))>((4'd10)!==(3'd2)))!=(((5'd26)&&(-3'sd1))<<((2'd3)<<(3'd6))));
  localparam [4:0] p13 = (^{1{(^{3{{1{(4'd0)}}}})}});
  localparam [5:0] p14 = (!(~&(|(!(((-5'sd0)&&(4'sd0))!==(&(2'sd0)))))));
  localparam signed [3:0] p15 = {(2'd2),(5'd13),(5'd7)};
  localparam signed [4:0] p16 = (3'sd1);
  localparam signed [5:0] p17 = (4'd6);

  assign y0 = ((~&(-(b4-a0)))?((|a0)>(~&a1)):(4'sd4));
  assign y1 = (((~(b3===b0))>=((b4==p2)==(p7==p7)))-(|(|((p11<<p5)/p10))));
  assign y2 = (+(4'd9));
  assign y3 = (p13+p7);
  assign y4 = (({3{p5}}>(p0))?((p12^p2)^~(p15-p12)):($unsigned(p8)&{p12,p2}));
  assign y5 = $signed((~|(((-(&{$unsigned({p13}),(a3^~p16)}))|({(~&{(p7?p4:p5)}),{a2,p1,a5}})))));
  assign y6 = (((-b0))/a3);
  assign y7 = ((~&b1)===(&b2));
  assign y8 = (({{2{a4}}}>{(-b0),{3{b2}}})!=={{3{b5}},{3{b0}},(a5&a1)});
  assign y9 = (p5<<<p3);
  assign y10 = (^(^(~|(+((p7==b0)-(^p9))))));
  assign y11 = ((~|p2)>>(a2-p5));
  assign y12 = ((|(&(~^(~&p8))))?(~&$signed((|(-p0)))):$unsigned((~^(~^(p11)))));
  assign y13 = (({{b2,p8},$unsigned(a0)}==((p15?a3:b3)|(^p7)))<(^{{b2,a0},(p6?b0:a0),{{b1}}}));
  assign y14 = (((p12^a0)<={b1,b1})>=(2'd3));
  assign y15 = (&({2{p7}}?{3{p9}}:(6'd2 * p12)));
  assign y16 = (2'sd1);
  assign y17 = (((-b3)?(^b5):(b0>=b3))?(|(~|(|(b1?a2:b1)))):((b5?b5:a1)?(a2&a3):(b4?a5:a5)));
endmodule
