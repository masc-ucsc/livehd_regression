module expression_00946(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(5'd22));
  localparam [4:0] p1 = (~|{2{{3{(4'd4)}}}});
  localparam [5:0] p2 = (((-5'sd12)<<(2'sd0))?((-2'sd1)>(-3'sd2)):{2{(5'd26)}});
  localparam signed [3:0] p3 = (({(2'd3)}?((3'd6)&&(5'd5)):(4'd3))?{((5'd13)+(-3'sd1)),(-(5'd22)),((2'd3)>>(3'd0))}:(|(~{(3'd7),(-5'sd0),(3'd0)})));
  localparam signed [4:0] p4 = {(~(5'sd3)),((3'sd0)?(-2'sd1):(-5'sd1)),(~|(-4'sd0))};
  localparam signed [5:0] p5 = (((^((-2'sd0)|(2'd3)))>{((3'd4)?(5'd19):(2'd1))})!=(((-5'sd8)!==(5'd29))?((2'd0)>(5'd22)):(|(2'd0))));
  localparam [3:0] p6 = {{({(-5'sd6),(5'sd8)}<<{((3'sd0)!==(3'd5))}),(((5'sd15)===(5'd27))<<<((5'sd14)|(-2'sd1)))}};
  localparam [4:0] p7 = (~^{3{{4{(3'd5)}}}});
  localparam [5:0] p8 = (5'd26);
  localparam signed [3:0] p9 = (~((~&(+{(5'sd6),(-5'sd4)}))&(((4'sd1)<(-3'sd1))+((4'd14)!=(-3'sd0)))));
  localparam signed [4:0] p10 = ((5'd22)!==(5'd1));
  localparam signed [5:0] p11 = ((((3'd5)>>(5'sd8))-((5'd17)>=(-3'sd1)))<=(((4'd9)===(4'd0))==((3'sd1)^(2'd3))));
  localparam [3:0] p12 = {((2'd3)>=(2'd0)),((4'd8)>>>(3'd2))};
  localparam [4:0] p13 = (&((((3'sd2)?(2'd0):(3'd3))!=((4'sd3)>>(5'd11)))|(((3'sd2)<=(3'sd3))==(4'd2))));
  localparam [5:0] p14 = {3{(|(4'd8))}};
  localparam signed [3:0] p15 = (~&((+(-5'sd12))^(3'd4)));
  localparam signed [4:0] p16 = (!(2'd1));
  localparam signed [5:0] p17 = ((((-3'sd3)==(4'd0))^~((5'd14)^~(3'd5)))|(((-3'sd1)^~(5'sd15))^~((2'd0)-(3'sd0))));

  assign y0 = ((p1?p15:p8)?{(~^(~^p11))}:{3{p1}});
  assign y1 = (|(&p14));
  assign y2 = (({b0}?(p7?p1:a3):(p6?a4:a1))?((p1?a0:p7)?(p13?p6:p16):{p0}):({a3,p6,p9}?{p12}:{p12}));
  assign y3 = (((2'd0)<=(&p8))!=((p12!=p12)<<{4{a2}}));
  assign y4 = ((&b3)===(-3'sd1));
  assign y5 = (((p4>a3)<<$unsigned((b5<<<p2)))<<$signed(((6'd2 * a0)>>(p7<p6))));
  assign y6 = (~^(~(5'd2 * (4'd2))));
  assign y7 = {2{{1{$signed({2{(b4?p5:a5)}})}}}};
  assign y8 = {{{p3,p14},{p6,p13},(p1?p14:b5)},((p12&&p2)?{p13,b1,p9}:(a1?b3:a2))};
  assign y9 = {{3{{b2,p4,p7}}},({{2{p3}},(p6>a3)}+((p9^b0)&{b0,a2}))};
  assign y10 = (^(~|(2'd0)));
  assign y11 = {{b5,p17}};
  assign y12 = (((b3<<a3))^(a4^~a1));
  assign y13 = (((a3===a2)<(5'd2 * p7))?((a0|a1)<={2{p0}}):((a3!=p2)>>(p12+a5)));
  assign y14 = {2{(&{1{({{b1,b3}}-(p10?p6:p8))}})}};
  assign y15 = {1{{{1{(~^(~|{(a1===a5)}))}},{4{(-a2)}},({2{b4}}>>(~(~^p12)))}}};
  assign y16 = ({1{((a4<<b1)|(6'd2 * a1))}}&{4{p1}});
  assign y17 = ({3{a1}}?(~&a4):{2{p15}});
endmodule
