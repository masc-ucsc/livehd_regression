module expression_00461(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(((2'd1)?(4'd13):(3'd2))?((-5'sd1)>=(-5'sd10)):{(3'd5)}));
  localparam [4:0] p1 = ((((2'd1)-(3'd3))>>((-3'sd2)-(2'd2)))!=(((5'd25)>(-2'sd0))<<{(3'd0),(-4'sd0),(5'sd3)}));
  localparam [5:0] p2 = {4{((3'sd3)?(4'd9):(3'd5))}};
  localparam signed [3:0] p3 = ((^((3'd0)?(4'd5):(5'd1)))==(((-3'sd2)?(-5'sd10):(-3'sd0))!=((5'd29)?(-3'sd1):(4'sd4))));
  localparam signed [4:0] p4 = (2'sd0);
  localparam signed [5:0] p5 = (~^(-((2'd3)!==(&((5'd6)||(-4'sd7))))));
  localparam [3:0] p6 = ({4{(~(4'd1))}}!={1{{3{(~^(-5'sd10))}}}});
  localparam [4:0] p7 = (5'd12);
  localparam [5:0] p8 = {(~(&(+(~&{((5'sd1)&&(5'd29)),(4'sd7)}))))};
  localparam signed [3:0] p9 = (4'sd6);
  localparam signed [4:0] p10 = ((((3'd1)>=(2'd3))==={(5'd25),(5'sd3),(-3'sd1)})-(~|{(4'd14),(4'd2)}));
  localparam signed [5:0] p11 = ((5'd10)?(~(~^{4{(5'd30)}})):{4{(2'd1)}});
  localparam [3:0] p12 = {4{{3{(-3'sd2)}}}};
  localparam [4:0] p13 = ((2'd1)|(&{1{((!(2'sd1))+((5'd4)>>(3'd2)))}}));
  localparam [5:0] p14 = (((-3'sd2)?(2'sd0):(2'd0))?{4{(2'sd1)}}:((3'sd0)>>>(3'sd3)));
  localparam signed [3:0] p15 = ((((3'd6)>>(-3'sd1))>((2'd0)&&(2'd2)))<(((2'd1)<=(-5'sd10))>(^(-3'sd1))));
  localparam signed [4:0] p16 = (((5'sd13)?(2'd3):(4'sd2))-((2'd1)?(2'd0):(-3'sd2)));
  localparam signed [5:0] p17 = (~&{((-2'sd1)<<<(4'sd5)),((5'sd8)>>(2'sd0))});

  assign y0 = {b2,b4};
  assign y1 = ({2{(b5?b0:b0)}}>=((~&{2{b3}})?(!(b5^a2)):$unsigned((+b4))));
  assign y2 = (({3{(p9<=p6)}}>>({3{p9}}>{1{p12}}))&&(^((^(~&{3{a3}}))<({3{p17}}<<(a1&b0)))));
  assign y3 = ((p5?b3:a4)?(|(a1?b2:b4)):(b2?b1:b4));
  assign y4 = {1{{1{{1{(!{3{{3{(|b3)}}}})}}}}}};
  assign y5 = (~^((p11<=p6)>=(b5==b2)));
  assign y6 = (((p4!=p1)?(!{p13,p8}):(~|(p8?p16:p9)))<=(~|(((a1>>>a4)+(a0|b0))===(b2?b0:b4))));
  assign y7 = ((6'd2 * (p12^p6))>>>((p6&p16)));
  assign y8 = (6'd2 * (4'd2));
  assign y9 = (((p17?p7:p2)?(p8|b1):(a3?a4:b1))?((p17+b5)?(a3&&p16):(b2==p17)):((p13?b0:a2)>>(p5?p8:b5)));
  assign y10 = {b1,b5};
  assign y11 = (-{$signed($signed({2{((a1>>>p12)^~(4'd1))}})),{(^(p2-p16)),(p5<p5),(-4'sd5)}});
  assign y12 = ({2{p8}});
  assign y13 = $signed(a4);
  assign y14 = {3{{3{(p13?p17:p4)}}}};
  assign y15 = (b3?a0:a5);
  assign y16 = (2'd2);
  assign y17 = $unsigned({1{{1{(-((~&(|{p9,p0}))))}}}});
endmodule
