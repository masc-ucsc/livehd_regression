module expression_00053(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'd2)?(5'd26):(2'd1))?((-4'sd1)?(3'd7):(4'd10)):{((2'd1)?(2'sd0):(4'd11))});
  localparam [4:0] p1 = {2{(5'd2 * (3'd5))}};
  localparam [5:0] p2 = {2{(2'd2)}};
  localparam signed [3:0] p3 = {(2'd3),(-5'sd4),(5'd23)};
  localparam signed [4:0] p4 = ((-2'sd0)|{{((-3'sd0)+(-2'sd0))},((5'd13)?(4'sd6):(4'd0))});
  localparam signed [5:0] p5 = {2{{1{(((5'd19)===(2'sd1))&((3'sd3)>=(2'sd1)))}}}};
  localparam [3:0] p6 = (2'd1);
  localparam [4:0] p7 = (((~(5'd27))?(|(3'd2)):(!(4'd14)))?(((2'sd1)?(2'd0):(4'd0))?((-3'sd0)?(4'sd5):(3'sd0)):(~(-5'sd15))):((|(3'd3))?((-4'sd2)?(3'd7):(5'sd12)):((-3'sd3)?(3'd6):(-3'sd0))));
  localparam [5:0] p8 = (&{{{(-4'sd7),(3'd3)}},{2{(4'd7)}}});
  localparam signed [3:0] p9 = (+(+(-5'sd3)));
  localparam signed [4:0] p10 = {2{{4{{(3'sd0)}}}}};
  localparam signed [5:0] p11 = {4{(5'sd13)}};
  localparam [3:0] p12 = {3{{3{(4'd13)}}}};
  localparam [4:0] p13 = (((5'd21)>(3'd2))!==(2'd3));
  localparam [5:0] p14 = (4'd13);
  localparam signed [3:0] p15 = (|{(~&{3{((3'd6)?(-2'sd0):(-3'sd0))}})});
  localparam signed [4:0] p16 = {{3{(-5'sd3)}},{1{(-4'sd0)}},({1{(5'd17)}}<=((5'd15)?(4'd4):(3'sd2)))};
  localparam signed [5:0] p17 = ((5'd11)||(-5'sd3));

  assign y0 = (a3==a1);
  assign y1 = (|(-4'sd3));
  assign y2 = ((-4'sd2)?(a5!==a3):(3'd6));
  assign y3 = (4'd8);
  assign y4 = {({(b3>a5)}>>(b0<<a3))};
  assign y5 = $unsigned({2{p8}});
  assign y6 = $signed((((a4^~b4)!=(a2!==b5))>>(4'd2 * $unsigned(b3))));
  assign y7 = $unsigned((2'sd0));
  assign y8 = (4'sd3);
  assign y9 = $signed(((4'sd6)));
  assign y10 = ((^{{{(b4>=p13)}}})-(5'd23));
  assign y11 = {3{(b0<p11)}};
  assign y12 = (^((5'd11)?(p6?p16:p7):{3{p14}}));
  assign y13 = ((+(b3&&p7))==(!(^b2)));
  assign y14 = (~|((2'sd0)));
  assign y15 = (~^(-2'sd1));
  assign y16 = (2'd3);
  assign y17 = (|(~^(~{2{{4{{2{p9}}}}}})));
endmodule
