module expression_00668(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-4'sd2);
  localparam [4:0] p1 = ({3{((-2'sd0)!==(3'd0))}}-({3{(2'd1)}}<<(|{3{(2'd0)}})));
  localparam [5:0] p2 = (((-2'sd0)-(4'sd3))!==((-4'sd2)===(-3'sd0)));
  localparam signed [3:0] p3 = {4{((4'sd1)!=(5'd29))}};
  localparam signed [4:0] p4 = (4'sd2);
  localparam signed [5:0] p5 = ((((3'd7)?(5'sd1):(-5'sd5))>=(-5'sd7))>(((5'sd2)*(5'sd7))/(2'd0)));
  localparam [3:0] p6 = ((((4'd8)==(3'd2))?((5'd20)^~(5'sd15)):((2'd3)>>(2'd1)))|(((3'd3)==(4'sd6))>>>((3'sd1)?(5'd13):(3'd6))));
  localparam [4:0] p7 = ((((5'd0)&&(2'sd1))=={2{(5'd14)}})^(~|({2{(5'sd8)}}^((2'd1)<<(3'sd1)))));
  localparam [5:0] p8 = (&(~((((2'sd1)>=(-5'sd10))==((5'd15)^(3'd5)))!=(!({(2'd2),(5'd12),(-3'sd3)}+{(3'sd3),(4'd14)})))));
  localparam signed [3:0] p9 = (((5'sd3)?(2'd3):(-2'sd1))?{4{(3'd1)}}:((-5'sd7)===(-2'sd1)));
  localparam signed [4:0] p10 = ({(-2'sd1),(5'd0)}?((4'd0)?(4'd11):(-4'sd5)):{(-4'sd3),(-4'sd5)});
  localparam signed [5:0] p11 = ((((5'd20)<<(4'sd6))<<(+(~&(5'sd6))))|(~(~|((~|(2'sd1))!=={3{(3'd2)}}))));
  localparam [3:0] p12 = ((~&(+((-5'sd6)?(2'd2):(3'd4))))?(|((4'd10)?(3'd3):(2'd3))):(^((4'sd4)?(5'sd8):(5'd5))));
  localparam [4:0] p13 = {4{{(3'd2),(2'd0)}}};
  localparam [5:0] p14 = {3{(5'd8)}};
  localparam signed [3:0] p15 = (~|(+{((~(+{(3'sd3),(5'd4),(3'd2)}))&&{(!((-5'sd11)?(2'd3):(-5'sd14)))})}));
  localparam signed [4:0] p16 = {1{(4'd3)}};
  localparam signed [5:0] p17 = ((3'sd1)&(-3'sd1));

  assign y0 = (5'd8);
  assign y1 = ((~^((a5<<b5)<=(-(b3^~p9))))?(&($unsigned(a2)?(~a3):(a0))):$unsigned((~&($signed(a4)|$unsigned(p1)))));
  assign y2 = ((-3'sd3)!=(((6'd2 * p14)>=(p15<=p0))&(2'd2)));
  assign y3 = ((p4?p11:p10)?(p17<<p13):{2{b4}});
  assign y4 = ((3'sd0)?(~&(p15?p16:p0)):(2'sd1));
  assign y5 = (3'd2);
  assign y6 = ((((4'sd0)^{a3})===(4'd10))-((-3'sd2)||(5'd15)));
  assign y7 = ($unsigned($unsigned($unsigned($unsigned($unsigned($unsigned($unsigned(b5))))))));
  assign y8 = ($unsigned(($signed(a1)<<(p7>>>p10)))?(3'd1):$unsigned((-4'sd6)));
  assign y9 = $unsigned(((5'sd4)>>(5'd30)));
  assign y10 = (~^({1{$unsigned(p12)}}?(3'd3):{4{p17}}));
  assign y11 = {2{{(b1!==b0),{p12}}}};
  assign y12 = $unsigned((!(($signed(p1))/p9)));
  assign y13 = (4'd2 * $unsigned((p10?p8:p0)));
  assign y14 = (~^{(!(~^{p7,p9,a5})),{(~^{p12})},{b3,p10,a0}});
  assign y15 = ($unsigned({{1{a3}}})?(b2?b3:p4):({3{a5}}&&(6'd2 * b2)));
  assign y16 = ((p10>>p13)&{4{p11}});
  assign y17 = (&(5'sd14));
endmodule
