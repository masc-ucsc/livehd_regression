module expression_00663(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~{{(-3'sd2),(3'sd2),(5'd7)},(5'sd7),(4'd5)})||(~^(|(((-3'sd1)?(5'sd3):(-3'sd0))==((-3'sd0)?(4'd7):(5'sd8))))));
  localparam [4:0] p1 = (|((4'sd3)?(2'd1):(4'd12)));
  localparam [5:0] p2 = (!(5'd20));
  localparam signed [3:0] p3 = (!(~^(5'd16)));
  localparam signed [4:0] p4 = ({4{(3'd1)}}!=({4{(-2'sd1)}}!={2{(5'd5)}}));
  localparam signed [5:0] p5 = ((&((5'd28)?(-4'sd5):(4'd11)))?(~((-4'sd7)^(2'sd0))):((3'd3)?(3'sd3):(5'd25)));
  localparam [3:0] p6 = ((3'sd2)<<({3{(3'sd0)}}<<{(4'd6),(2'sd1)}));
  localparam [4:0] p7 = {4{((3'sd3)+(3'd1))}};
  localparam [5:0] p8 = (6'd2 * {1{((2'd0)|(3'd4))}});
  localparam signed [3:0] p9 = ({1{((2'd3)&&(-3'sd3))}}>{2{((-3'sd3)<=(5'd17))}});
  localparam signed [4:0] p10 = ((4'd11)>>>(4'sd1));
  localparam signed [5:0] p11 = (3'sd3);
  localparam [3:0] p12 = ((^(-2'sd1))&(-2'sd1));
  localparam [4:0] p13 = (((3'd0)+(2'd0))/(4'sd6));
  localparam [5:0] p14 = (((-3'sd1)>>(5'd11))>>>{(2'd3),(2'd1),(-2'sd0)});
  localparam signed [3:0] p15 = {(~|(5'sd14)),{(3'sd0),(-4'sd4)}};
  localparam signed [4:0] p16 = {((-5'sd6)?(3'sd2):(-5'sd7)),{3{(2'd2)}}};
  localparam signed [5:0] p17 = (~|(~^(+(^(~(~&((~^(2'sd1))*(3'd1))))))));

  assign y0 = (((~^a1)&(p6<<<p4))?((&a1)-(p3|p5)):({1{a4}}?(p3<<p1):(p2<<<p6)));
  assign y1 = (&((((b1||a4)<=(a4-a4))!==(~(a5^b4)))>((4'd2 * (+a1))>((~a4)==(^b3)))));
  assign y2 = ({1{{4{(3'd0)}}}}>>$unsigned((~&$unsigned(((3'd0)&&((a2-b1)))))));
  assign y3 = {2{{4{{2{p11}}}}}};
  assign y4 = $unsigned((($signed((5'd2 * p6))<=((|p12)/a3))<<<((b0?p2:a4)+((a4^~b4)+(p3!=a1)))));
  assign y5 = (((b3&&p9)>=(b4===b0))<<((p17<p9)>>(p0-a3)));
  assign y6 = ((!(~|(-a1)))?{1{(~(-2'sd1))}}:{4{a4}});
  assign y7 = ((((p14==p3)-(^b2))=={4{a5}})>>{4{(p17>>p10)}});
  assign y8 = {3{{(~{b3})}}};
  assign y9 = (!{4{((~b3)<<<(-p8))}});
  assign y10 = ((((b3?a5:a5)<<<(a0<<b4))!==(b5?b5:a0))<<(4'd15));
  assign y11 = {1{{{4{a4}},(b0+a2),{2{a2}}}}};
  assign y12 = {{4{a0}},(~^{b2,p6}),{(5'd2 * b2)}};
  assign y13 = (4'sd7);
  assign y14 = (2'd2);
  assign y15 = ($signed(((+p9)))&(5'd20));
  assign y16 = (~(5'sd13));
  assign y17 = ((5'sd4)==(5'd7));
endmodule
