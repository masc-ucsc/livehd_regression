module expression_00843(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(4'sd0));
  localparam [4:0] p1 = {1{(!{{{(2'sd1)},(|(3'sd0))},(&(~|(|(|(2'd2)))))})}};
  localparam [5:0] p2 = (-3'sd1);
  localparam signed [3:0] p3 = ((2'd0)>>>(4'sd7));
  localparam signed [4:0] p4 = (4'd7);
  localparam signed [5:0] p5 = {((5'sd10)<(-2'sd1)),(2'd0),{(3'd7),(2'd0),(4'd3)}};
  localparam [3:0] p6 = ((|(2'sd1))^(5'd2 * ((3'd4)!=(5'd9))));
  localparam [4:0] p7 = (((2'd1)<<(3'd4))>=((5'd13)<<<(-5'sd15)));
  localparam [5:0] p8 = ((4'd14)>>((3'd1)&&((4'd0)||(3'sd2))));
  localparam signed [3:0] p9 = (!{2{(4'd9)}});
  localparam signed [4:0] p10 = {(2'd3),(4'sd1)};
  localparam signed [5:0] p11 = (({(5'd18),(4'd7),(2'd1)}+((3'd3)==(-2'sd0)))-(((3'sd0)>>(5'd23))-((-4'sd0)?(2'd2):(5'd19))));
  localparam [3:0] p12 = {(((5'd5)!==(4'd4))&{4{(-3'sd1)}})};
  localparam [4:0] p13 = (((~{2{(5'd18)}})-{1{((5'sd8)>(3'd7))}})<<<((!((2'sd0)&&(4'sd0)))^((2'sd0)|(-4'sd7))));
  localparam [5:0] p14 = (4'd2 * ((2'd0)==(2'd1)));
  localparam signed [3:0] p15 = (((^(-2'sd1))?{(-4'sd2)}:(!(5'sd6)))?((+(-4'sd3))?{3{(4'd13)}}:{(5'd12),(-3'sd0),(3'd4)}):((-(5'd10))?{4{(4'sd0)}}:(|(-3'sd2))));
  localparam signed [4:0] p16 = (-((((-2'sd1)>(3'd7))-((3'sd0)<<<(-2'sd0)))&&(-(+((|(5'd6))^~((3'd2)|(-2'sd0)))))));
  localparam signed [5:0] p17 = (-3'sd0);

  assign y0 = {(b3>>>a3)};
  assign y1 = (|(^a5));
  assign y2 = ((-3'sd2)|(5'sd14));
  assign y3 = $unsigned(a4);
  assign y4 = (~&$unsigned({1{(5'sd1)}}));
  assign y5 = {{{{3{p5}}},{p2,p17}},({2{a1}}==(p1&&b1)),({3{p16}}<{p13,p16})};
  assign y6 = {2{{1{p11}}}};
  assign y7 = (5'd29);
  assign y8 = (!(~^(-(~&p13))));
  assign y9 = ((~|({2{{4{a3}}}}<=((~&p4)>={4{b3}})))^(((~&p7)<<<(~a4))<((a3==p4)&(+a5))));
  assign y10 = (4'd7);
  assign y11 = ((-(p7<=p10))^(p12-p17));
  assign y12 = (4'd3);
  assign y13 = (|p17);
  assign y14 = (((a2)?$unsigned(b0):{4{b2}})>>($unsigned({4{p4}})));
  assign y15 = (4'sd3);
  assign y16 = (~|((~(^p1))|(p2|a1)));
  assign y17 = (4'd2 * (p0<=p13));
endmodule
