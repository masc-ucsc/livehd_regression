module expression_00306(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~((3'sd3)>>{1{(+(4'd11))}}));
  localparam [4:0] p1 = (((2'd2)<<(5'sd6))|(&(-(5'sd3))));
  localparam [5:0] p2 = (^({2{((2'd2)==(3'd4))}}&&{3{(-2'sd1)}}));
  localparam signed [3:0] p3 = {(~^{(3'd6),(2'd1),(-3'sd3)}),(^{(-(5'sd4)),(4'sd0)}),(~^(2'd1))};
  localparam signed [4:0] p4 = (3'sd0);
  localparam signed [5:0] p5 = ((~^(2'sd0))?(2'sd0):{1{((4'sd3)==(3'd4))}});
  localparam [3:0] p6 = (3'sd2);
  localparam [4:0] p7 = (-4'sd1);
  localparam [5:0] p8 = ((((4'd6)!=(-5'sd1))||((4'sd3)<(5'sd14)))-((5'sd3)?(-5'sd15):(4'd4)));
  localparam signed [3:0] p9 = (((-4'sd2)!=(-5'sd12))===(~&(|(2'd3))));
  localparam signed [4:0] p10 = (~(+(((+(-3'sd0))^~(2'sd0))<{2{(4'd2)}})));
  localparam signed [5:0] p11 = ({{3{(2'sd0)}},{2{(5'sd2)}},((-3'sd3)?(2'd0):(5'd25))}?{{(-3'sd3),(2'd1),(3'd1)},(~&(2'd1)),((4'd3)>=(2'sd1))}:(((5'd13)?(5'sd1):(-2'sd0))<<(~|(2'd0))));
  localparam [3:0] p12 = ((((-5'sd15)!=(2'd1))==(6'd2 * (4'd15)))!=(((5'd27)<<<(4'sd0))<{1{((5'd28)>>(3'd1))}}));
  localparam [4:0] p13 = (+(+((~((-3'sd3)|(2'd2)))!=(~((3'd4)===(3'd5))))));
  localparam [5:0] p14 = ({4{(3'd6)}}?((4'sd2)?(-2'sd1):(2'd2)):(4'd9));
  localparam signed [3:0] p15 = {2{{2{((5'sd8)>>>(-5'sd0))}}}};
  localparam signed [4:0] p16 = (2'sd0);
  localparam signed [5:0] p17 = ((2'd1)?(((-5'sd14)>>(2'd0))^~(6'd2 * (5'd3))):{(^(3'd0)),((4'd12)<<(4'sd6))});

  assign y0 = (~^(-(~{(-(a5^~p15)),(3'd0)})));
  assign y1 = ({4{p10}}?{{p4,p5},{p2,p2},{p10,p6,b3}}:(~^{1{{4{p10}}}}));
  assign y2 = ((4'sd6)?{p0,a4,b0}:{p6,b4});
  assign y3 = ((+{b5,p1,p6})-$signed(((~|p7))));
  assign y4 = (({{b3,p16,p7}}||(4'd6))||(((|a4)>{3{b5}})==={3{a0}}));
  assign y5 = (((a3&&a4)>>{2{p16}})?((4'sd4)>=(2'sd1)):(~|{4{b4}}));
  assign y6 = (+((a0|b5)?{p0,p7,b2}:{$signed(p1)}));
  assign y7 = (2'd1);
  assign y8 = (^(({4{p7}}?(p7&p4):(a0?p14:a4))&((!(a1>=b0))?(p7|a0):{2{p11}})));
  assign y9 = {1{(~|{2{(~^(~&{2{b0}}))}})}};
  assign y10 = ((~|$unsigned((-5'sd11)))?({4{b3}}?(b3?b5:a5):(^a4)):(-5'sd15));
  assign y11 = ((a0>=b1)==={a5,a4,b1});
  assign y12 = (4'sd6);
  assign y13 = {1{(($signed({2{b3}})&&((b5&b1)))!==((+(~|a4))>=$unsigned({4{b2}})))}};
  assign y14 = $signed(((4'd2 * b1)?(p2):(-2'sd0)));
  assign y15 = ({4{(a5?b2:b5)}}!==$unsigned({1{((a4==b5)?(a1<<<a5):(b1?a0:b5))}}));
  assign y16 = (($signed(a4)+{b4,a1})^((b1<a4)>>(b5&a4)));
  assign y17 = (-3'sd0);
endmodule
