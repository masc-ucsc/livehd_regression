module expression_00792(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(!(2'sd0)));
  localparam [4:0] p1 = {4{{3{(4'd0)}}}};
  localparam [5:0] p2 = (+{4{(~((-4'sd2)&&(-2'sd1)))}});
  localparam signed [3:0] p3 = {4{(3'd2)}};
  localparam signed [4:0] p4 = (~^{(-5'sd8),(2'd1)});
  localparam signed [5:0] p5 = ((|((5'd21)?(4'sd3):(3'sd1)))!==((3'd4)|((-5'sd8)>(-4'sd7))));
  localparam [3:0] p6 = ({(-2'sd0)}?(!(3'sd1)):(+(2'd3)));
  localparam [4:0] p7 = {1{{{(+(-3'sd3))},{1{(~&(4'd9))}},{(-2'sd1),(2'd2),(4'd10)}}}};
  localparam [5:0] p8 = ((((4'sd3)<=(-4'sd4))===((3'sd0)|(3'd2)))&(((4'd13)?(2'd1):(-4'sd3))>>(-4'sd7)));
  localparam signed [3:0] p9 = (((5'sd8)^(2'd2))<<((-3'sd3)&&(-3'sd3)));
  localparam signed [4:0] p10 = {4{(3'd1)}};
  localparam signed [5:0] p11 = (~(3'sd3));
  localparam [3:0] p12 = ((3'sd2)>=(2'd1));
  localparam [4:0] p13 = (~^(((5'd0)/(3'd1))<=((4'd2 * (4'd12))<<((4'sd7)||(4'd15)))));
  localparam [5:0] p14 = {2{{(5'd9),(3'd7)}}};
  localparam signed [3:0] p15 = ({3{(&(2'd0))}}||(((5'd29)^(2'd3))?((3'sd1)?(3'd4):(5'sd3)):{2{(2'sd1)}}));
  localparam signed [4:0] p16 = (~^(-(~|((&(^((4'd1)?(4'd3):(2'd3))))?((-4'sd4)?(5'd18):(3'd2)):(~&((-3'sd0)?(3'd2):(4'd1)))))));
  localparam signed [5:0] p17 = {{4{(3'd0)}},{1{{2{(-4'sd5)}}}}};

  assign y0 = ((-(2'd3))>=(-4'sd0));
  assign y1 = ((~((~a4)^$unsigned(p0)))?$unsigned(((^a3)-(&a4))):((p6*b4)==(!p10)));
  assign y2 = {{3{{1{(p7||p16)}}}},({3{((p6))}})};
  assign y3 = {((b1!==a5)===(a4>>>b0)),((|(~|p2))<<(a5===a1)),(3'd2)};
  assign y4 = ({{b4,a4,b5},{a4,b2,a1}}+(4'd12));
  assign y5 = $signed({{(3'sd1)}});
  assign y6 = {$unsigned({2{$signed($unsigned(p14))}})};
  assign y7 = (b1>>a5);
  assign y8 = (({4{p13}}^(4'd2))?(3'sd2):((-5'sd0)>>>(b5+p1)));
  assign y9 = (a3?a4:p10);
  assign y10 = {(({1{b1}}?(b3<=a5):(-4'sd7))),(3'd2),{1{(^(a5?a3:a4))}}};
  assign y11 = (((+p3)>(p14<<<p11))>>((p11)<=$signed(p3)));
  assign y12 = (p10==a0);
  assign y13 = $signed((((p7?p15:p1)&&$unsigned({1{(p1<=p16)}}))));
  assign y14 = ((b2|b3)%b4);
  assign y15 = ((p13?p10:p0)*(b5^~b4));
  assign y16 = (|$signed(((~^$unsigned((!p7)))!=(&(+(!a3))))));
  assign y17 = {2{(((b0>>>b1)>(a0===b4))<((~p14)<<<(b1>a3)))}};
endmodule
