module expression_00924(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{{2{{(2'sd0),(4'd7),(3'sd2)}}}}};
  localparam [4:0] p1 = (2'd1);
  localparam [5:0] p2 = (!((4'd1)<<<(5'd2)));
  localparam signed [3:0] p3 = ({(5'd24),(-2'sd1)}>=(~^(2'sd1)));
  localparam signed [4:0] p4 = (~&{3{(-{1{(4'd4)}})}});
  localparam signed [5:0] p5 = (~^((5'd11)>>(4'd12)));
  localparam [3:0] p6 = ((+((-2'sd1)?(2'd2):(-3'sd3)))?({3{(5'd3)}}?((5'd6)?(2'sd1):(3'd7)):((-4'sd4)||(3'sd3))):(~({2{(4'd3)}}!=(|(3'd7)))));
  localparam [4:0] p7 = {4{(!(3'd1))}};
  localparam [5:0] p8 = (((4'sd0)?(3'sd0):(3'd5))||{4{(3'd7)}});
  localparam signed [3:0] p9 = (^((|(2'd0))^~(~|(3'sd0))));
  localparam signed [4:0] p10 = (((-3'sd1)>=(3'd2))!==(5'd2 * (2'd3)));
  localparam signed [5:0] p11 = {3{((5'd13)^(-3'sd0))}};
  localparam [3:0] p12 = (((3'd4)?(5'd25):(4'd9))<(+(4'd11)));
  localparam [4:0] p13 = (&((~&{4{(-5'sd0)}})<{1{(2'd0)}}));
  localparam [5:0] p14 = ({(3'sd3),(3'd2),(5'sd11)}===((4'd14)?(2'd0):(-4'sd7)));
  localparam signed [3:0] p15 = ((-5'sd2)==(2'd3));
  localparam signed [4:0] p16 = ((+(6'd2 * (|(5'd21))))-{4{(2'd2)}});
  localparam signed [5:0] p17 = (!{{(^{{(~|(4'd10))}}),{{(4'sd3)}},{(~(3'sd1))}}});

  assign y0 = {(((b5||p3)?(b0<<<b0):(4'd2 * p7))),((a0?b2:a3)?(p10>=p16):{p12,p9,a2})};
  assign y1 = ((~^a0)?(3'd1):(a0?a4:a3));
  assign y2 = (4'd2 * {p2,p8});
  assign y3 = ((a2^p13)|{3{p9}});
  assign y4 = ((5'd2 * p12)?$signed((a3+a4)):(p5?b4:p9));
  assign y5 = (-4'sd2);
  assign y6 = {4{p8}};
  assign y7 = {4{{{b5,b0,b1},(+a3),(^a3)}}};
  assign y8 = ((5'sd8)==(b0));
  assign y9 = (+(~(3'd0)));
  assign y10 = $unsigned({2{({p13,b4}>(p6-a3))}});
  assign y11 = {3{(~&((~&p11)==(a2&&b5)))}};
  assign y12 = (5'd3);
  assign y13 = ((-{2{((6'd2 * a1)>=(b0===a1))}})||(~|(!((b0!==a5)<<<{1{(a4&a5)}}))));
  assign y14 = (3'sd3);
  assign y15 = (b4^~p15);
  assign y16 = (b3*b4);
  assign y17 = ((5'sd5));
endmodule
