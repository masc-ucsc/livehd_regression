module expression_00734(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^(-4'sd5));
  localparam [4:0] p1 = ({2{(-3'sd3)}}<={2{(-5'sd10)}});
  localparam [5:0] p2 = ((^(3'sd1))?(~&(2'sd0)):((5'd18)>>>(4'd12)));
  localparam signed [3:0] p3 = (((((4'd7)>=(5'd6))<((5'd5)<(3'd2)))==(((4'sd0)^(4'd13))|((-2'sd0)+(5'sd3))))|((((2'd3)<<(5'd27))/(5'd29))&(((-3'sd0)/(2'd2))!=((5'sd12)!=(5'd8)))));
  localparam signed [4:0] p4 = (!(((!(5'd29))?((4'd8)^~(3'sd3)):((3'd7)==(5'd2)))^~(~^((4'sd3)?(4'd12):(4'd8)))));
  localparam signed [5:0] p5 = (&((!((&((4'd6)^(4'd10)))>((5'd25)<<<(-2'sd0))))^((-(^(4'sd0)))!==((-5'sd4)<(2'sd1)))));
  localparam [3:0] p6 = (^(5'd15));
  localparam [4:0] p7 = (~^(~((-5'sd2)^~(~&(-4'sd6)))));
  localparam [5:0] p8 = (~(4'd13));
  localparam signed [3:0] p9 = (((3'sd0)+(5'd3))+(5'd4));
  localparam signed [4:0] p10 = (!((3'sd3)<<(((-2'sd1)-(3'd7))!=((-3'sd3)<<<(4'sd7)))));
  localparam signed [5:0] p11 = (!(4'd12));
  localparam [3:0] p12 = ((-2'sd0)&((3'sd1)?(-4'sd4):(4'd9)));
  localparam [4:0] p13 = (-5'sd11);
  localparam [5:0] p14 = {1{{1{({2{{2{(-4'sd0)}}}}?(((-3'sd2)?(-5'sd10):(-5'sd13))?((5'd14)?(5'sd1):(5'd3)):((2'd0)?(-4'sd2):(2'd1))):{4{(2'd1)}})}}}};
  localparam signed [3:0] p15 = {2{{2{{4{(5'd28)}}}}}};
  localparam signed [4:0] p16 = {{{{(5'd18)},{(-4'sd2),(4'd10)},(+(5'sd8))}}};
  localparam signed [5:0] p17 = ((4'd11)?(3'd3):(4'sd4));

  assign y0 = (~|{(!{3{(~^{4{b5}})}})});
  assign y1 = (~&(~^$signed((!(~&(|(b0>>b3)))))));
  assign y2 = (({b2}!==(|a4))>>(~^(4'd2 * {3{b2}})));
  assign y3 = (|($unsigned((~|(a4>=a3)))>=(a5?b0:b4)));
  assign y4 = (-2'sd1);
  assign y5 = {3{$signed({1{(p9>>b2)}})}};
  assign y6 = (~^({p0,a2,p5}?(~^(a1?a4:b0)):(|{3{p3}})));
  assign y7 = ($unsigned((3'sd2))?$signed(((5'd23))):$unsigned($unsigned((3'sd2))));
  assign y8 = ((b3!==a5)!==$unsigned($signed(a1)));
  assign y9 = (b2^p15);
  assign y10 = (|({(a1||p8),{a2,p12,p5}}<<(3'd5)));
  assign y11 = (~&(b5?b5:p9));
  assign y12 = $signed((2'd2));
  assign y13 = ({1{{2{(-3'sd1)}}}}>>>(-4'sd2));
  assign y14 = ($signed({$unsigned(p1),(~^p4)}));
  assign y15 = {{b1,p9,p17},{b1,b4,p15},$unsigned(b1)};
  assign y16 = ((~{2{(p15||p11)}})?((5'd9)^{1{(p10|p9)}}):((b1?p8:b1)>(p5<<p0)));
  assign y17 = (~|(((a2)?(~^b0):(~&a5))?((~|(~|$unsigned(b0)))):(-(!(p15?b5:a3)))));
endmodule
