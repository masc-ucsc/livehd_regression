module expression_00686(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(5'd9),(3'sd2),(4'd4)},{3{(2'd1)}}};
  localparam [4:0] p1 = {1{{{3{(3'd7)}},{(5'd10)},{4{(5'sd11)}}}}};
  localparam [5:0] p2 = {3{(!{3{(3'd3)}})}};
  localparam signed [3:0] p3 = ((~^((-2'sd1)+((3'd7)&(4'sd2))))&&(((3'd7)?(2'd3):(3'sd3))?((3'd0)?(3'd5):(2'd0)):{3{(3'd4)}}));
  localparam signed [4:0] p4 = {4{((3'd3)?(2'sd0):(5'd7))}};
  localparam signed [5:0] p5 = (|((~&(~&((-3'sd2)|(2'd0))))>(+(((3'd0)^~(2'sd0))>((2'd1)<<<(5'd1))))));
  localparam [3:0] p6 = (6'd2 * ((4'd7)?(5'd7):(5'd11)));
  localparam [4:0] p7 = {1{{({2{{(3'd7)}}}?(((2'sd1)?(2'd0):(4'sd2))=={(4'sd3),(-5'sd0),(5'd8)}):(((5'sd9)?(5'd1):(2'd3))|{3{(2'sd1)}}))}}};
  localparam [5:0] p8 = ((3'sd0)?(~&(~^(2'd2))):(-3'sd1));
  localparam signed [3:0] p9 = (!(~&(~^((!(5'd6))-(~|(-5'sd4))))));
  localparam signed [4:0] p10 = (&(&((4'sd5)?(3'sd2):(2'd3))));
  localparam signed [5:0] p11 = (2'd1);
  localparam [3:0] p12 = {2{((2'd0)?(-3'sd2):(-5'sd14))}};
  localparam [4:0] p13 = ((+(((3'd6)!=(2'd2))<(~|((2'sd0)+(-5'sd4)))))>>>{1{(~^{2{(!((-5'sd11)===(2'sd1)))}})}});
  localparam [5:0] p14 = ({1{{1{{1{{2{{1{(3'd1)}}}}}}}}}}!=={{3{(5'd1)}},{(5'd25),(-5'sd13)}});
  localparam signed [3:0] p15 = ({{1{(3'sd1)}},((3'sd1)!==(4'd13))}!=={{(-2'sd0),(4'sd2)},{(3'd0),(-4'sd3),(5'd12)}});
  localparam signed [4:0] p16 = ((6'd2 * {4{(2'd0)}})?{1{(((2'sd0)?(-4'sd3):(-3'sd0))<<((3'sd0)>(-5'sd5)))}}:(+({2{(2'd2)}}!==(^(3'd3)))));
  localparam signed [5:0] p17 = (5'sd14);

  assign y0 = $unsigned(($signed((2'd0))));
  assign y1 = {4{$signed((2'd3))}};
  assign y2 = (|(|(~&p0)));
  assign y3 = $signed((~$unsigned((~&($unsigned((5'd1))?$unsigned((3'sd2)):(a0?a5:a4))))));
  assign y4 = {1{{1{({(^b0),$unsigned(b1)}=={2{(b2!==b4)}})}}}};
  assign y5 = ((|(!(-4'sd1)))?(-{(4'd2 * p6),(+b4),{3{b0}}}):({1{(a1===b4)}}!==(-5'sd15)));
  assign y6 = (~|((b1&&p13)+(~&b0)));
  assign y7 = (3'd0);
  assign y8 = (p14?p0:p14);
  assign y9 = $signed($unsigned((3'd2)));
  assign y10 = {$unsigned(((-(b0<=b3))>>>((b1<<b0)))),(({a3,a2,p17}>>>{b3,b4})&(|((a1))))};
  assign y11 = (2'd2);
  assign y12 = (~&(p5|p11));
  assign y13 = (~|a4);
  assign y14 = {{1{(6'd2 * {3{a2}})}}};
  assign y15 = {({(a0>>b1)}&{(a4<b5),(p6>a3)}),{({b4,p15}||(p12+p2))}};
  assign y16 = (~|{4{(p3?a3:p15)}});
  assign y17 = (((-({2{a2}}<$unsigned(p7))))>=(~|{4{a1}}));
endmodule
