module expression_00614(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((5'sd13)==(-3'sd0))>((3'd0)>>>(2'd1)))+(-((~|(3'd4))-(-2'sd0))));
  localparam [4:0] p1 = {((4'sd6)?(2'd1):(4'd2)),{1{(~|{(-4'sd0),(5'sd2),(4'sd2)})}}};
  localparam [5:0] p2 = (((3'd3)?(3'd7):(4'd13))?((-3'sd3)%(2'd3)):((2'd0)-(-2'sd0)));
  localparam signed [3:0] p3 = (({(2'd2),(3'd3)}&(~|{(2'd0)}))<=(+{2{{2{(-3'sd3)}}}}));
  localparam signed [4:0] p4 = (((5'd23)&&(3'sd0))?(~&((3'sd0)?(-3'sd1):(5'd8))):((2'sd0)?(2'd0):(-2'sd0)));
  localparam signed [5:0] p5 = {((4'd3)<<(2'sd0)),(&(-5'sd9)),(&(3'd7))};
  localparam [3:0] p6 = (!(~^(~^{((5'd29)?(4'sd6):(3'd4)),{(-4'sd7),(3'd6),(4'd14)},{(-3'sd1),(2'd0),(-5'sd15)}})));
  localparam [4:0] p7 = (((5'd21)+(5'd15))?((2'd3)?(4'sd4):(-3'sd1)):{3{(5'd10)}});
  localparam [5:0] p8 = (4'd0);
  localparam signed [3:0] p9 = (~&({2{(+(4'sd6))}}<={2{{4{(4'd12)}}}}));
  localparam signed [4:0] p10 = (!((2'd0)!==(5'd12)));
  localparam signed [5:0] p11 = {(3'd4),(4'sd1),(-2'sd1)};
  localparam [3:0] p12 = (5'd28);
  localparam [4:0] p13 = (^(-3'sd2));
  localparam [5:0] p14 = (!(-4'sd7));
  localparam signed [3:0] p15 = (5'd16);
  localparam signed [4:0] p16 = {2{(((3'd5)>(5'd19))&&{1{(4'd10)}})}};
  localparam signed [5:0] p17 = ((5'sd4)?(5'sd10):(3'sd1));

  assign y0 = {$unsigned((|{{p2,p8,p16},(-5'sd14)}))};
  assign y1 = $unsigned({{{p1,p11,p7},(|{p13,p2}),(!{3{p0}})},(5'd9)});
  assign y2 = (&(4'sd4));
  assign y3 = (((($signed(p5))==(p11?p15:p2)))?((p3<<<p1)!=(p12?p16:p4)):((p12?p17:p12)<<<$signed((p3?p10:p16))));
  assign y4 = {2{{p5,b4,p10}}};
  assign y5 = ((p7?p15:p17)?(p14?p1:p3):((p7<=p15)<<(p13-p11)));
  assign y6 = (&{3{(|p3)}});
  assign y7 = {({$unsigned({{p11,p14,p7},(b2>b0)})}>$signed((2'sd1)))};
  assign y8 = (-4'sd2);
  assign y9 = ((~^(p16?p0:p9))?((a3||a5)===(b4>=b5)):({p14,p9,b0}?(p17<<p0):(p13!=p5)));
  assign y10 = (((a5&b5)%a5)<<<$signed($signed($signed((p7-b0)))));
  assign y11 = ($unsigned(($unsigned($signed(p3))<<{4{p0}}))-(4'd2 * {2{p13}}));
  assign y12 = $signed((!$signed((+$signed($signed(p8))))));
  assign y13 = {{2{((p10?p13:b2)?(p3?a1:a1):{a4,b1,p9})}}};
  assign y14 = (-3'sd0);
  assign y15 = (4'sd2);
  assign y16 = (~^$signed((p6?p9:p2)));
  assign y17 = {3{$signed(({3{b1}}<<(b2!==a3)))}};
endmodule
