module expression_00263(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(-5'sd8)};
  localparam [4:0] p1 = (^(3'd2));
  localparam [5:0] p2 = {(^((-3'sd1)>>(4'sd4))),(~&{(-5'sd9),(2'd3)}),({2{(4'sd2)}}!==((3'd2)<<(3'd2)))};
  localparam signed [3:0] p3 = (4'sd7);
  localparam signed [4:0] p4 = (((-4'sd7)?(4'd5):(-5'sd15))?(~&(!(5'd19))):((3'd7)?(3'd4):(4'sd5)));
  localparam signed [5:0] p5 = (2'sd1);
  localparam [3:0] p6 = ({({(-3'sd2)}|((-5'sd7)&&(2'sd1)))}<<{((2'sd0)-(5'd13)),((4'd15)>>>(5'd8)),(-(2'sd0))});
  localparam [4:0] p7 = (-(2'sd1));
  localparam [5:0] p8 = ((5'd2 * ((4'd4)===(5'd23)))+(((2'sd1)*(2'sd0))!==((5'sd6)>>(2'd1))));
  localparam signed [3:0] p9 = ((4'd3)/(3'd3));
  localparam signed [4:0] p10 = (^(((5'sd11)>(4'd3))?(~(-2'sd1)):{4{(2'd1)}}));
  localparam signed [5:0] p11 = ((2'd0)?(2'd2):(-3'sd2));
  localparam [3:0] p12 = (((4'd2)?(3'sd1):(4'd11))===(!(2'sd1)));
  localparam [4:0] p13 = (~|(2'd3));
  localparam [5:0] p14 = {(4'd14),(-2'sd0),(-2'sd0)};
  localparam signed [3:0] p15 = (5'd26);
  localparam signed [4:0] p16 = ({1{(5'sd1)}}?((-5'sd9)||(-5'sd11)):((-5'sd6)^~(-4'sd0)));
  localparam signed [5:0] p17 = ((!((4'd14)+(-2'sd0)))?{((4'd5)-(3'd4)),((-3'sd1)<<(2'd0))}:({(4'sd7),(-5'sd15),(4'd10)}!=((5'sd15)?(5'd23):(4'd2))));

  assign y0 = ((-4'sd0)>>>({a1,a5}<<<(a0||b5)));
  assign y1 = (((~|(a1<<p14))?(b4>>a3):{a2,a1})^~(~^((a5<<a4)?(b1==b1):(a0?b2:a5))));
  assign y2 = (~(~^(((-p2))?(|$unsigned(p10)):{(p9?p8:p13)})));
  assign y3 = (5'sd6);
  assign y4 = ($signed((b3<a0))!==($unsigned(b4)>{1{a1}}));
  assign y5 = {1{(+(({3{{3{b3}}}}?{4{p17}}:((b0?p5:b2)!=(a3>p17)))))}};
  assign y6 = ({4{(p5>>a0)}}&(~(^((b3+b4)<<<(~|a4)))));
  assign y7 = {(^((b3>a2)?(p8?p1:p11):(b2?p16:b3)))};
  assign y8 = (p16?b4:p1);
  assign y9 = (4'd5);
  assign y10 = (p3|p1);
  assign y11 = ({a3,p10,p12}^((p7+b5)^~(p11<=p0)));
  assign y12 = (((~|(p17?b2:a2))^~{3{(b2?a4:p1)}})&&(({1{p15}}?{2{a2}}:(a2?b2:b3))==(5'sd5)));
  assign y13 = (((5'd14)?{b2}:{a5,p5,b3})?{(5'd31),{1{a5}},{b1,b2}}:(!(+(a5?a5:a1))));
  assign y14 = {b0,p12,p4};
  assign y15 = ((p4?p6:b5)?(b5?a2:p0):(p6^~a4));
  assign y16 = ({2{b2}}&(b3?p6:a3));
  assign y17 = {{{{p17,b5}},{{p13,p15,a5},{p7,p15}},{{p14,p16}}}};
endmodule
