module expression_00434(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{3{(-5'sd2)}}}};
  localparam [4:0] p1 = (~|((~((4'sd2)>>((4'd1)?(4'd13):(5'd31))))!=(3'd2)));
  localparam [5:0] p2 = {2{((5'd30)+(3'sd0))}};
  localparam signed [3:0] p3 = (+(~&{{4{((3'd7)?(-2'sd1):(5'd4))}}}));
  localparam signed [4:0] p4 = {{1{(!((5'sd6)?(4'd0):(-3'sd3)))}},{{(-5'sd6),(4'sd7),(2'sd1)}}};
  localparam signed [5:0] p5 = (4'd8);
  localparam [3:0] p6 = ((~|((5'd17)^(3'sd2)))>>>((4'sd2)?(4'd15):(5'd16)));
  localparam [4:0] p7 = (((3'sd2)>((-2'sd1)==(2'sd1)))>(((2'sd1)^~(3'd3))^{1{((3'd3)>(3'd3))}}));
  localparam [5:0] p8 = (|(6'd2 * (&{1{(3'd5)}})));
  localparam signed [3:0] p9 = ((((2'sd0)&(2'd0))|((5'sd13)>>(5'sd9)))!==((|((-4'sd5)<<(-2'sd0)))||(+((-5'sd6)!=(2'd3)))));
  localparam signed [4:0] p10 = ((-3'sd0)+(-4'sd0));
  localparam signed [5:0] p11 = (((3'd2)||(2'sd1))<=((5'sd13)+(3'd1)));
  localparam [3:0] p12 = (((4'd4)|(3'd5))>((5'd1)<(5'sd5)));
  localparam [4:0] p13 = ((3'sd0)||(2'sd1));
  localparam [5:0] p14 = ((+(~^(3'd3)))/(4'd10));
  localparam signed [3:0] p15 = ((~(-3'sd2))?((4'd2)?(-3'sd3):(3'd5)):{(4'sd3),(2'd0),(-5'sd11)});
  localparam signed [4:0] p16 = {(-3'sd0),(~&(~|(!(2'd2)))),((5'd4)?(-3'sd0):(-2'sd1))};
  localparam signed [5:0] p17 = ((-3'sd1)?(4'sd5):(4'd0));

  assign y0 = {4{(4'd2 * (3'd0))}};
  assign y1 = ((b2<=a3)!=(p5<p12));
  assign y2 = ((b1-p16)<(^p9));
  assign y3 = ((~((p8<<b1)<=(a5-a2)))^~(2'sd0));
  assign y4 = (&(~^(-((p15&p9)<<(&p11)))));
  assign y5 = (-2'sd1);
  assign y6 = $unsigned((-((^(+({2{b4}}<<<(~(-a0)))))<<<($unsigned((^(p9?a3:b2)))||(p10?p14:a4)))));
  assign y7 = {(~{2{p12}}),(!(~^p5)),(p1^~p2)};
  assign y8 = ({(p4+p17),(p2|p0),(p7)}&((p5-p0)?(p10?p3:p9):(p8?p11:p13)));
  assign y9 = (((~|b1)+(b0^~b0))>>((~^b5)===(a1-b2)));
  assign y10 = (-4'sd7);
  assign y11 = (^(&(|($signed(((~^$unsigned(p5))|((3'd1))))>>>($signed((+(~a4)))===$signed((~^(a2^~a5))))))));
  assign y12 = (~^(((b1?b2:a2)===({b1,b3}-(b0)))&&(5'd26)));
  assign y13 = ({{(&(p11<<p7))},($unsigned(p9)-(^b2))}<<<((&(~|(a3-p4)))-{1{((|p10)>>{4{p10}})}}));
  assign y14 = (-3'sd1);
  assign y15 = (($signed(p17)?(p0?p0:b4):$signed(a2))?($signed(a1)?$unsigned(b5):$unsigned(p11)):((p6?p17:p4)?$signed(p3):(a1?p7:a5)));
  assign y16 = ((2'sd0));
  assign y17 = ((4'd6)>{a0,p6,b1});
endmodule
