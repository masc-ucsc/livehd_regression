module expression_00911(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(&((5'd24)>=(2'd0)))}};
  localparam [4:0] p1 = ((5'd2 * {2{(5'd17)}})>={1{(((4'd5)+(-5'sd3))^(6'd2 * (3'd3)))}});
  localparam [5:0] p2 = (~^((~&(~((-2'sd1)<<<(3'd6))))>>{(-(5'd14)),((-5'sd15)<=(-5'sd7))}));
  localparam signed [3:0] p3 = (5'd2 * (^(~(4'd13))));
  localparam signed [4:0] p4 = ((((3'd2)?(2'd2):(2'sd0))?((-4'sd1)>(3'd3)):(5'sd0))||(~&(-3'sd1)));
  localparam signed [5:0] p5 = (((^(+(|(2'sd0))))-(-((2'd3)===(-4'sd4))))!==((&((3'd7)^(-4'sd1)))===(-((-2'sd1)===(-4'sd0)))));
  localparam [3:0] p6 = (~&((2'd1)|(2'd2)));
  localparam [4:0] p7 = ((&(5'd17))?(!(3'd7)):((-3'sd3)?(4'd11):(-5'sd9)));
  localparam [5:0] p8 = ((((-5'sd12)?(3'd7):(3'd6))+(~&(2'sd0)))?(((3'sd1)?(2'd1):(-2'sd0))>((3'd6)?(2'sd1):(-5'sd6))):((~(-4'sd5))+((2'sd0)==(5'd25))));
  localparam signed [3:0] p9 = {4{{3{(3'sd1)}}}};
  localparam signed [4:0] p10 = (|(2'sd1));
  localparam signed [5:0] p11 = ((((3'd7)>>>(-4'sd2))>((5'd31)<<<(2'd1)))>(~&((-4'sd2)<<(-5'sd15))));
  localparam [3:0] p12 = ((^(2'd1))^~{2{(3'd7)}});
  localparam [4:0] p13 = ((~|(4'sd1))<{4{(5'sd2)}});
  localparam [5:0] p14 = {2{(~&{(~(~&(~{3{(3'd7)}})))})}};
  localparam signed [3:0] p15 = (+((-(((4'd8)+(2'sd1))-((4'sd2)&(3'd3))))>>(!(~(((3'd6)===(4'd14))&&((3'sd3)<=(4'd9)))))));
  localparam signed [4:0] p16 = ((-(!(2'd0)))==(3'sd2));
  localparam signed [5:0] p17 = {2{(|(-(~^{1{(5'd7)}})))}};

  assign y0 = ((a3<=a5)&&(p8?p2:b3));
  assign y1 = $signed($signed((!(~{3{(~&{3{b0}})}}))));
  assign y2 = (((p17&&p0)<(~|p1))&(^((a3?p1:p4)||(p14|p13))));
  assign y3 = (((p16>>>b0)<{p11,p1,p7})!=(^((a0>p14)&&{2{a2}})));
  assign y4 = ((((p6<p5)&&{b1,p11})+{p0,a2,a3})&&{2{((5'd2 * b2)&(a0?a2:p9))}});
  assign y5 = {(b1),{p7},$signed(p6)};
  assign y6 = (~(+(^(((a2<<a1)!=(-5'sd5))<=(-5'sd5)))));
  assign y7 = {{p3,p12},{p16,p4},{p14,p16}};
  assign y8 = {3{$signed((~^(&a2)))}};
  assign y9 = (4'sd7);
  assign y10 = (({1{a5}}<={3{b4}})>>>((a4>=b1)&&{2{b5}}));
  assign y11 = ({1{((p3>>>p17)^(3'd1))}}>>>(2'sd1));
  assign y12 = $unsigned({$signed((!(($signed(({3{b3}})))<<{{(5'd11)}})))});
  assign y13 = $unsigned({((b3^~b4)?(a2):(a4?a2:p3)),{(^(^(a1?a1:b0)))}});
  assign y14 = ((~^$signed(b3))!={p17,b5,b3});
  assign y15 = ((a5==p7)^~(4'sd7));
  assign y16 = (b2>>>p9);
  assign y17 = (2'd2);
endmodule
