module expression_00049(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'd2)?(5'sd6):(-3'sd0))<(~((3'd4)^(4'd12))));
  localparam [4:0] p1 = ((+(|(!((-5'sd1)&&(3'sd3)))))>(!(5'd2 * ((4'd9)!==(5'd6)))));
  localparam [5:0] p2 = (~|(|(|(&(+(-2'sd0))))));
  localparam signed [3:0] p3 = (~|{(~((-5'sd12)-(2'd2))),{{(2'd3),(-4'sd0)}}});
  localparam signed [4:0] p4 = {(((4'sd1)&&(-2'sd0))!==((2'sd1)>=(-5'sd1))),{((2'sd1)^~(3'd6)),((2'sd1)<(4'sd6)),((4'd8)-(5'sd7))}};
  localparam signed [5:0] p5 = (+(({1{(2'd0)}}^~((-5'sd6)+(2'd3)))||(((3'd0)>>(4'sd7))!==((4'd11)&(2'sd1)))));
  localparam [3:0] p6 = {2{((3'd7)===(3'd2))}};
  localparam [4:0] p7 = (4'sd5);
  localparam [5:0] p8 = ((((4'd4)===(4'sd1))<=(~|(-3'sd1)))>>>(6'd2 * (&(3'd5))));
  localparam signed [3:0] p9 = ((&((3'd1)?(3'd2):(4'd7)))!==((4'sd1)?(5'd17):(-4'sd3)));
  localparam signed [4:0] p10 = (&(6'd2 * (~&((5'd25)?(2'd1):(2'd3)))));
  localparam signed [5:0] p11 = {{{(4'd9)},(~&(-5'sd2)),((2'sd0)?(-3'sd3):(4'd6))},{{(-2'sd1)},(~(5'd25))},(^{(4'd8),(2'd2),(3'sd0)})};
  localparam [3:0] p12 = ((4'sd7)!=(4'sd6));
  localparam [4:0] p13 = (({2{(-3'sd1)}}<=(6'd2 * (3'd1)))<<<(((4'sd1)<<(-5'sd7))&(~|(4'sd4))));
  localparam [5:0] p14 = (^(~&(2'd0)));
  localparam signed [3:0] p15 = {2{(6'd2 * ((3'd5)^(2'd2)))}};
  localparam signed [4:0] p16 = (((2'd1)>>(2'd0))?(!(+(3'sd0))):((2'd1)?(5'sd7):(3'sd1)));
  localparam signed [5:0] p17 = (&(~^(^((+(2'sd0))/(4'd4)))));

  assign y0 = ($signed((~&(~&{p10,a4})))?{(&p15),(b3===a0)}:($unsigned(a3)=={a1}));
  assign y1 = (((~&(a1|b4))^~(!(~^b0)))>((a5?b5:p4)?(~&a4):(b1?p13:b2)));
  assign y2 = $unsigned(((4'sd1)));
  assign y3 = (2'sd0);
  assign y4 = (!{2{({{3{p8}},(a3&&p14)}&&(&{3{p12}}))}});
  assign y5 = (&{2{((p2<<<p9)>>(~&(p13>p1)))}});
  assign y6 = (|((p3?p15:p16)?((a2?b4:b0)||{a4,p6}):(~(p3?a3:p13))));
  assign y7 = $signed({3{p13}});
  assign y8 = (~|(~&((!(a5>b2))&(4'd2 * b2))));
  assign y9 = {1{(b4?a2:b1)}};
  assign y10 = (!(^$unsigned($unsigned((3'd1)))));
  assign y11 = (~&({4{a0}}?(!b4):(4'd8)));
  assign y12 = ({3{(p6+p0)}}?((p17?p16:p9)?(p2&&p3):(p15<<<p16)):((!p11)<<{3{p1}}));
  assign y13 = (((p14+a1)||(b0>=a3))>>>{(p5<=p10),(2'd0),{b0,b0}});
  assign y14 = ((~&b0)>>(b3!=b1));
  assign y15 = (~^{2{({1{((b0^a4)^(a3-a4))}}==(-({1{a1}}^~{4{b3}})))}});
  assign y16 = {((a5?a1:b5)?(a0?a5:a4):(a1?p11:b0)),((p12?a3:b0)?{a2,b0,a4}:{b5,a0})};
  assign y17 = {1{$signed(({2{{1{(-5'sd14)}}}}))}};
endmodule
