module expression_00509(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd14);
  localparam [4:0] p1 = {(3'sd0),(2'd3),(4'sd5)};
  localparam [5:0] p2 = (((5'sd15)==(2'sd0))>>>((-3'sd3)!=(-5'sd3)));
  localparam signed [3:0] p3 = (|((-3'sd1)&(2'd1)));
  localparam signed [4:0] p4 = (4'sd7);
  localparam signed [5:0] p5 = (5'sd12);
  localparam [3:0] p6 = (&(!((-3'sd3)?(3'd6):(2'sd1))));
  localparam [4:0] p7 = ((~&(3'sd2))<<(4'd6));
  localparam [5:0] p8 = ((((4'd13)?(3'd5):(4'd4))||((3'd1)?(-2'sd0):(5'd10)))?((2'd0)?(2'd0):(4'd2)):((2'd3)<(6'd2 * (2'd3))));
  localparam signed [3:0] p9 = ((2'd1)-(4'd5));
  localparam signed [4:0] p10 = (!{{((4'd7)?(-4'sd1):(-3'sd0)),((5'd4)==(4'd15)),(~|(2'sd1))},((+(-5'sd5))?((-2'sd1)?(2'd2):(3'd4)):(4'd3)),(-4'sd3)});
  localparam signed [5:0] p11 = {4{{2{(4'd1)}}}};
  localparam [3:0] p12 = {1{((5'd0)?(3'sd3):(2'sd1))}};
  localparam [4:0] p13 = {{(3'd6)},((4'd2)&&(^((2'sd1)?(4'd14):(3'd1))))};
  localparam [5:0] p14 = ((((4'd13)?(5'd28):(4'sd7))!==(((3'd3)?(-5'sd2):(2'd0))|((3'd2)?(-2'sd1):(2'sd1))))+(((4'd1)&&(3'd7))?{((-4'sd0)?(4'd14):(4'd7))}:{1{((2'd1)?(3'd7):(2'sd1))}}));
  localparam signed [3:0] p15 = (-(-({(5'd10),(4'd2),(2'd1)}>(~(4'd3)))));
  localparam signed [4:0] p16 = (6'd2 * (-{3{(3'd3)}}));
  localparam signed [5:0] p17 = (5'd12);

  assign y0 = {{{((^(b2&&p5))>>((p6-p8)<(~^a0)))},(~^({p11,p7,p9}>(-{p11,p0})))}};
  assign y1 = (~&(~|{(-{{{a5,p15}}}),(&{{a1,p7,p0}}),(|(~^{a2,a2,a3}))}));
  assign y2 = (((p4?p13:a5)&(p8!=p8))^~{1{(!(|p13))}});
  assign y3 = ((&((!(b0==p15))/b4))+((4'd6)!=(~&(|(2'd1)))));
  assign y4 = {3{(^a4)}};
  assign y5 = {$signed({1{(2'd3)}})};
  assign y6 = ((-4'sd6)||((4'd2 * b1)|(+(a2||a4))));
  assign y7 = $unsigned((~|(((+(-3'sd0))?(5'sd12):(5'sd10)))));
  assign y8 = {3{{(a1-p14),{4{p16}}}}};
  assign y9 = (-4'sd5);
  assign y10 = ({3{b3}}?(~|(a5!=b2)):(b3?b5:a4));
  assign y11 = ((^((p14||p5)>{4{p3}}))<<(5'd13));
  assign y12 = {3{(|(&{2{(&a3)}}))}};
  assign y13 = {4{{a4,b2}}};
  assign y14 = (-((~|((|(a3?b3:p15))<{3{b5}}))>>>{1{(+{1{(2'd3)}})}}));
  assign y15 = {(p6?p11:b4),(p12?b1:p6)};
  assign y16 = (~^(a5?p6:b4));
  assign y17 = ((p6%p0)<<<(+(|p0)));
endmodule
