module expression_00806(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd2)<<<(-4'sd2))>=((2'd3)?(-3'sd3):(5'sd0)))?{4{(3'd6)}}:((4'd5)?(-2'sd0):(5'd8)));
  localparam [4:0] p1 = (((2'sd0)==(4'd13))>>((5'd14)&(3'd1)));
  localparam [5:0] p2 = ((-2'sd0)+(3'sd0));
  localparam signed [3:0] p3 = ((-3'sd3)%(-5'sd15));
  localparam signed [4:0] p4 = (({(-4'sd7),(4'd15),(2'd1)}>>((-2'sd1)!==(5'd0)))^~({(4'd4),(-2'sd1),(2'sd1)}>=((4'd11)<<(-2'sd1))));
  localparam signed [5:0] p5 = ({((4'd6)<<(2'd1)),{(5'd2),(2'sd1)},{(5'sd2),(4'd15),(3'd4)}}>={{{(4'sd1),(2'sd0)},{(-2'sd0)}},(((3'd0)>>(4'd7))==((4'd12)+(4'sd2)))});
  localparam [3:0] p6 = ({2{((4'sd1)||(5'd7))}}>>{1{{4{(2'd0)}}}});
  localparam [4:0] p7 = {((4'd4)?(3'd0):(2'sd1)),((3'sd0)?(2'd3):(-4'sd2))};
  localparam [5:0] p8 = (((-2'sd1)?(5'sd9):(-4'sd1))?(~^(~&((5'd26)?(3'd0):(3'sd1)))):(^((-3'sd3)?(3'd0):(5'd18))));
  localparam signed [3:0] p9 = ((~|(!((3'sd0)%(2'd1))))==(((5'sd6)+(-3'sd0))|((3'sd3)>=(-5'sd10))));
  localparam signed [4:0] p10 = ((&((5'd29)?(2'd0):(-3'sd0)))>>>((4'd4)&(-4'sd4)));
  localparam signed [5:0] p11 = (+{(4'sd7),(4'd13),(4'd15)});
  localparam [3:0] p12 = {1{{1{(5'sd4)}}}};
  localparam [4:0] p13 = (~^(~^((|((~(-2'sd0))&&(~^(3'd1))))!==(((2'd1)&&(5'd24))&(~^(-(2'd3)))))));
  localparam [5:0] p14 = ((((4'd0)?(5'd1):(3'd3))?{(3'sd0),(-5'sd10),(4'sd2)}:{(4'sd6),(-3'sd2)})?(((2'sd1)>>(-5'sd4))?{(2'd3),(2'd0)}:{(2'd2),(2'd2)}):(-2'sd1));
  localparam signed [3:0] p15 = ({2{((-3'sd0)+(4'd5))}}^(((5'd23)||(4'sd4))|((-5'sd11)<<(3'd4))));
  localparam signed [4:0] p16 = ((~((3'd1)||(2'd3)))?(6'd2 * ((5'd20)%(4'd7))):(-((3'd6)|(5'd26))));
  localparam signed [5:0] p17 = (((5'd14)>>((5'd17)?(-4'sd2):(-2'sd0)))^~(2'd1));

  assign y0 = (~|(~(~&(!({1{{2{b1}}}}?(~^{p3,a2,p7}):(~^(+(p1|p11))))))));
  assign y1 = (~|(b4&b1));
  assign y2 = $signed((|{2{{((a2>p7)),(p12?p3:p0)}}}));
  assign y3 = (b3<=p1);
  assign y4 = ((~|(~|(~{p17})))&$signed((5'd2 * (p0<<p7))));
  assign y5 = {{a4,b5,a4},{p17,b4},{(b3&p13)}};
  assign y6 = (-((-(!(4'd7)))^~{(5'd26),(~|((5'd14)!==(b3>>b0)))}));
  assign y7 = (-(4'd14));
  assign y8 = (((p4?p10:p8)-(p13>>>p10))>>>(3'sd2));
  assign y9 = (a5==b4);
  assign y10 = ((b0)!={4{b2}});
  assign y11 = {3{{3{a3}}}};
  assign y12 = ({2{{p5,p3}}}==(~($signed({p10,p2,b5}))));
  assign y13 = {({(+(~p8)),{2{p12}}}^~((({4{b5}}===(!a3)))))};
  assign y14 = (~&(a2<<p1));
  assign y15 = (((p5+p9)^~(p6/p4))<<((p14-p10)<=(p14>>>p17)));
  assign y16 = (~|((a0===b2)-(^p15)));
  assign y17 = (-((~^{b4,b5})?(|(!b4)):(-(-p8))));
endmodule
