module expression_00187(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&{3{((5'd3)+(-2'sd1))}});
  localparam [4:0] p1 = {3{(-5'sd1)}};
  localparam [5:0] p2 = ({1{((-4'sd2)?(3'sd3):(2'sd1))}}>=(|(((2'd1)+(3'd1))|(+(2'sd1)))));
  localparam signed [3:0] p3 = (-2'sd1);
  localparam signed [4:0] p4 = {(|(-2'sd1)),((2'sd1)&(5'd14))};
  localparam signed [5:0] p5 = (6'd2 * (3'd0));
  localparam [3:0] p6 = {4{(4'sd7)}};
  localparam [4:0] p7 = (&(~(-(((~^(-2'sd0))>(+(-5'sd7)))?(&(!(|(2'sd0)))):((^(-5'sd12))<((4'd7)?(4'd7):(3'd7)))))));
  localparam [5:0] p8 = {{(-2'sd0),(3'd7)},(4'd2 * (3'd0))};
  localparam signed [3:0] p9 = ({(-3'sd3),(2'd0)}&(5'd28));
  localparam signed [4:0] p10 = (~^{(2'sd0),((^(3'd3))!={(-5'sd12)}),(4'd4)});
  localparam signed [5:0] p11 = (5'd4);
  localparam [3:0] p12 = ((2'sd1)&(3'd3));
  localparam [4:0] p13 = (-2'sd0);
  localparam [5:0] p14 = {3{((-3'sd0)?(5'sd3):(2'd1))}};
  localparam signed [3:0] p15 = ((5'd17)?(2'd1):(3'sd2));
  localparam signed [4:0] p16 = (4'sd2);
  localparam signed [5:0] p17 = {4{((3'd6)|(4'sd4))}};

  assign y0 = (-4'sd1);
  assign y1 = $signed((((b1!==b4)>=(^(^p8)))));
  assign y2 = (({2{p14}}|{p16,p16})&&(^{1{(p14<p14)}}));
  assign y3 = {((a3>a5)<=(+p1)),$unsigned(((-5'sd7)||$signed(a0))),(-3'sd1)};
  assign y4 = (-(((a4+p1)?(p1>>p10):(!a2))?((a5?b3:b0)!==(~a1)):((a1?b2:a0)>>(&b3))));
  assign y5 = (4'd1);
  assign y6 = {1{{2{({2{a2}}?(4'sd7):(3'd6))}}}};
  assign y7 = ({(p2-p16),{p6,p17}}?{1{(^{(p11^~p11)})}}:((p11>>>p11)|(p17^p1)));
  assign y8 = (((a5===b2)==(p9-a4)));
  assign y9 = $unsigned((({3{p3}}^~(~(~|p10)))!=({3{p4}}>>>(p6^~p14))));
  assign y10 = (3'd5);
  assign y11 = (((a2==p5)||{p16,p5})>>>{1{{a5,p4,b2}}});
  assign y12 = {$unsigned((3'd3))};
  assign y13 = {4{{4{p13}}}};
  assign y14 = (((~^(((b0!=a2))===(-4'sd2))))>>>(~&((p14?p7:p1)&&(~^(p9?p7:p5)))));
  assign y15 = {1{((p13!=p0)^{4{p17}})}};
  assign y16 = (^{1{(-5'sd0)}});
  assign y17 = $signed(({1{(({2{a1}})&(~^(b1)))}}-($unsigned({4{p2}})<<<({1{b1}}^(b2<b5)))));
endmodule
