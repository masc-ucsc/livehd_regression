module expression_00948(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^((2'sd0)>>>(-5'sd11)))>>>{(4'd3),(2'd1),(5'd26)});
  localparam [4:0] p1 = (2'd2);
  localparam [5:0] p2 = ((((3'd5)%(5'sd15))*((-5'sd1)<<(3'sd1)))>>>(((5'd23)<(5'sd1))?((2'd3)-(3'sd0)):((-5'sd6)>>(-5'sd8))));
  localparam signed [3:0] p3 = {{{1{(5'sd4)}},{3{(4'sd2)}}},{4{(4'd10)}},{(4'sd2),(4'sd6),(4'd10)}};
  localparam signed [4:0] p4 = {{{{(-3'sd0)},((5'd0)|(2'd3))},(^((3'sd1)?(2'sd1):(2'sd1))),((2'd1)?(2'sd1):(-2'sd1))}};
  localparam signed [5:0] p5 = {(4'd0)};
  localparam [3:0] p6 = {3{(|(2'd2))}};
  localparam [4:0] p7 = {2{(^{4{(3'd7)}})}};
  localparam [5:0] p8 = ((~^(~^(~(~&((-5'sd1)&(3'd0))))))^~(~^((!(^(5'sd10)))^((5'sd1)/(2'sd0)))));
  localparam signed [3:0] p9 = (+((-(+(((2'd3)<<<(3'sd2))*((-5'sd4)>=(2'd3)))))-(((3'd2)>>>(-2'sd1))<((4'd4)<<(5'sd2)))));
  localparam signed [4:0] p10 = (!((~&((5'sd0)<(2'sd1)))?((2'd0)?(4'sd4):(2'd0)):((-5'sd2)?(-4'sd6):(-2'sd1))));
  localparam signed [5:0] p11 = (((2'd3)>>>(2'd0))?((3'sd2)?(2'd3):(2'd2)):(&(4'd0)));
  localparam [3:0] p12 = ((&(((5'd9)||(2'sd1))>=(-4'sd5)))>=(~{4{{1{(-4'sd6)}}}}));
  localparam [4:0] p13 = ((((4'd7)>(-5'sd2))<=(|(2'd2)))&&((~^(-5'sd6))==(|(4'd3))));
  localparam [5:0] p14 = {4{(4'd0)}};
  localparam signed [3:0] p15 = (^(+(~{2{(4'sd2)}})));
  localparam signed [4:0] p16 = ((~^((4'sd4)?(-5'sd5):(5'sd9)))?(~|(((2'sd1)?(-3'sd2):(5'd2))!=(-(5'd2)))):((-(2'sd1))^((3'd4)%(5'd23))));
  localparam signed [5:0] p17 = (&{4{(-2'sd1)}});

  assign y0 = $signed({b0,b2,a1});
  assign y1 = (|$signed({2{{2{{a4,a1,a3}}}}}));
  assign y2 = ((|{3{$signed(b4)}})<<<$signed({3{$signed(b1)}}));
  assign y3 = (3'sd3);
  assign y4 = ((p1?b0:p16)/p1);
  assign y5 = {{(~^(!(!{(5'd7)})))}};
  assign y6 = (~|p0);
  assign y7 = (|((5'd2 * (&(b0%b1)))-(~|(4'd2 * (5'd13)))));
  assign y8 = (-3'sd1);
  assign y9 = {3{{b4,b0,b2}}};
  assign y10 = (a2?a0:b4);
  assign y11 = (|(+(~^((p8||p7)%p10))));
  assign y12 = (((a3<a1)<<(p15||p0))^~((b5===a4)^~(-p2)));
  assign y13 = ((a2^a1)<<(a3?a1:b0));
  assign y14 = ((-{{4{(~|p10)}}})-(&(({2{a3}})===((a3>>b3)===(a0>>>a0)))));
  assign y15 = {{{2{p5}},{2{p16}},(b0>=p14)},{(p5?p3:p6)},{{p13},(p8?p8:p11),(p9>p6)}};
  assign y16 = {4{(($unsigned((p1?a1:a0))))}};
  assign y17 = (|(((b3?p13:p2)>>(!p7))<{2{(p1?p8:p3)}}));
endmodule
