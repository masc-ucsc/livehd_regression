module expression_00391(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(~&(&{1{{{2{(2'sd0)}},(3'sd0),(~(&(4'd12)))}}}))};
  localparam [4:0] p1 = (3'sd1);
  localparam [5:0] p2 = (((-4'sd0)?(4'd2):(2'd0))?(~^(^((-5'sd10)?(5'd11):(-5'sd9)))):((4'd15)?(5'd18):(4'sd0)));
  localparam signed [3:0] p3 = (~|((~(~(3'd1)))<<(&{(4'sd6),(2'd0)})));
  localparam signed [4:0] p4 = {2{((+(3'sd0))?((-5'sd1)<<(-3'sd3)):(^(2'd3)))}};
  localparam signed [5:0] p5 = {3{(3'd4)}};
  localparam [3:0] p6 = {{{(4'd9),(4'd8)},{(5'sd13),(5'd30),(-5'sd2)}},{{(-5'sd1),(-3'sd1),(-4'sd5)},{(4'd5),(2'sd0),(2'd1)}}};
  localparam [4:0] p7 = {(+{((3'd0)!=(4'sd4)),((-2'sd0)|(4'd10))}),(((-4'sd5)&(2'sd0))&&{(4'd1),(-2'sd0)})};
  localparam [5:0] p8 = {1{(-(-5'sd12))}};
  localparam signed [3:0] p9 = (-4'sd5);
  localparam signed [4:0] p10 = ({(2'sd1),(-3'sd0),(5'd10)}<((4'sd0)?(2'd0):(-4'sd7)));
  localparam signed [5:0] p11 = ({4{(3'sd2)}}?({3{(4'd14)}}?(-(2'd2)):{2{(-4'sd6)}}):(|(~|{3{(5'sd2)}})));
  localparam [3:0] p12 = {{(4'sd1),(-3'sd3)}};
  localparam [4:0] p13 = (((3'd6)^(-3'sd2))*((2'sd1)<<<(5'd1)));
  localparam [5:0] p14 = ((5'sd4)?(-2'sd1):(2'sd1));
  localparam signed [3:0] p15 = ((+((-5'sd12)?(-2'sd1):(4'sd7)))?(((5'd16)?(-3'sd2):(5'sd3))|{(3'sd1),(-3'sd0),(5'd13)}):(&{(5'd31),(3'sd2)}));
  localparam signed [4:0] p16 = (3'd7);
  localparam signed [5:0] p17 = ((2'd3)<<<(4'd9));

  assign y0 = (((p12?p7:p4)||(p3?p15:p3))?{(p13?p9:p13)}:((a1^~p11)&&(p16?p5:p15)));
  assign y1 = ({3{(b3>p17)}}||({a4}-(p6^a4)));
  assign y2 = (((5'd20)^(-5'sd14))<$unsigned({4{(b1||b2)}}));
  assign y3 = (4'd2 * (6'd2 * p14));
  assign y4 = ((4'd0)^{1{{1{(2'd3)}}}});
  assign y5 = (-$unsigned((~^(&(~(a4<a2))))));
  assign y6 = ((&(((p7<<<p4)*(p16<=p6)))));
  assign y7 = ((-3'sd2)+((-2'sd0)^(~^(p4^p11))));
  assign y8 = ((p15^p5)?{2{a1}}:(p10^~p16));
  assign y9 = (((b5?p15:p11)?(2'd2):{4{p8}})-(+(5'd17)));
  assign y10 = (p8?p14:p4);
  assign y11 = ((^(p13>>p7))?(~{{p14}}):((p7?p15:p13)^~(-p1)));
  assign y12 = (|(a0===b3));
  assign y13 = ({1{(b5===a4)}}?{1{{p4,a0,a1}}}:{(a1>=b2)});
  assign y14 = (~((b3?a2:a4)/b1));
  assign y15 = ($signed((a4&&a4))==={1{((2'sd1))}});
  assign y16 = (3'd6);
  assign y17 = {2{(-5'sd14)}};
endmodule
