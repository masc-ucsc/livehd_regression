module expression_00450(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(4'd8));
  localparam [4:0] p1 = ((^(4'd5))?((5'd2)?(-2'sd0):(3'd3)):(-(-5'sd4)));
  localparam [5:0] p2 = (~^(~|(~&{((-(-5'sd0))==={(4'sd0),(5'd19)}),{4{(2'sd1)}},{4{(5'd19)}}})));
  localparam signed [3:0] p3 = (~^(~^(-(&(|{1{(&{4{(-2'sd1)}})}})))));
  localparam signed [4:0] p4 = (((2'd3)==(-4'sd2))/(5'sd10));
  localparam signed [5:0] p5 = ((2'd2)+(4'sd3));
  localparam [3:0] p6 = ((((3'd4)?(2'd3):(4'd15))>=((2'sd1)?(4'sd5):(5'd24)))!==(~^(((4'd10)===(4'd6))!=((-2'sd0)?(3'd2):(-3'sd0)))));
  localparam [4:0] p7 = {3{(2'd2)}};
  localparam [5:0] p8 = ((&(5'd2 * (4'd10)))<={(-4'sd2),(5'd18),(2'd2)});
  localparam signed [3:0] p9 = ({3{(-3'sd3)}}||(4'd2 * {1{(3'd2)}}));
  localparam signed [4:0] p10 = ({(((3'sd3)?(2'd1):(3'd3))>>((3'sd0)!==(2'sd0)))}<=(((5'sd14)?(5'd10):(5'sd6))<=((3'sd0)^(4'd9))));
  localparam signed [5:0] p11 = (((5'd21)<(2'sd0))^((2'd0)&(4'sd6)));
  localparam [3:0] p12 = ((~((3'd4)>=(-5'sd12)))?((5'sd12)?(4'd3):(5'd3)):(&((2'd3)?(2'sd1):(4'd5))));
  localparam [4:0] p13 = (4'sd4);
  localparam [5:0] p14 = {3{{(4'd14),(4'd7),(2'd3)}}};
  localparam signed [3:0] p15 = ((~|{4{((2'sd1)>>>(5'd2))}})==={(|(|(3'sd0))),(+(!(-2'sd1))),{(2'd3),(2'd1),(3'd2)}});
  localparam signed [4:0] p16 = ((4'sd6)>(4'd13));
  localparam signed [5:0] p17 = ((~(4'd11))*(~|(4'd14)));

  assign y0 = (((-(p8?a5:p0))>>>(p10+b0))<(~^{$unsigned(b0),(^a5),(b5^p6)}));
  assign y1 = {(4'd15),(!((&(p4-p1))-{p0,p3,p15}))};
  assign y2 = (({4{b4}}^~(a2||b2))!=((p10<=a0)==(a3>>>a2)));
  assign y3 = (((a2>>b2)^~(b2<<<b1))-(~&{4{(b5<<b5)}}));
  assign y4 = ((p0&&a1)||(b2?p17:p2));
  assign y5 = $signed((((5'd2 * a2)^(a2?b0:b3))!=(((b0-a1)===$unsigned((b1===a5))))));
  assign y6 = (!(~(((p8)-(a1?a2:a2))?(p2?p2:b4):{p7,p12,p11})));
  assign y7 = (!((^(a3>>a0))&&(b1>>>a0)));
  assign y8 = (((^(b5%b2))||(~^(b5%b4)))?((~(b5-b4))*(-(a2+b3))):(-(|((p8?b3:a4)<<(5'd2 * a1)))));
  assign y9 = ((a0?a2:b1)?$signed({(a1?b5:b3)}):{p17,a1,a0});
  assign y10 = (4'd8);
  assign y11 = (-2'sd0);
  assign y12 = $signed(($unsigned({2{(p14>>>b3)}})?$unsigned(((a0?b3:b0)?$signed(b0):$unsigned(a5))):((b0!==a2)!=$unsigned({1{p11}}))));
  assign y13 = (|{4{(-(~&{p14,a3}))}});
  assign y14 = ((~&b4)>>(b3?a5:a4));
  assign y15 = ((4'sd6)||((p9<<p3)<=(b2^~p5)));
  assign y16 = (+{2{{3{a3}}}});
  assign y17 = (((~|(a1>=p6))!={p1,p16,p0})^(-((!(p5-b4))|(p2^p12))));
endmodule
