module expression_00218(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(4'd3));
  localparam [4:0] p1 = ((-5'sd6)||(3'd0));
  localparam [5:0] p2 = (~(+({((2'd1)?(4'd10):(5'd4)),(~(3'd6))}<=(|({(4'sd5),(2'sd0),(4'sd3)}|{(2'd0),(2'sd1),(-3'sd0)})))));
  localparam signed [3:0] p3 = (3'd4);
  localparam signed [4:0] p4 = ((((3'd4)|(-3'sd3))&((5'd8)==(3'sd1)))!={{1{(-5'sd11)}},{3{(5'sd1)}},((3'd5)?(2'd1):(3'd6))});
  localparam signed [5:0] p5 = (6'd2 * (5'd12));
  localparam [3:0] p6 = (4'sd0);
  localparam [4:0] p7 = (|{(&(^{((5'd1)?(-5'sd8):(3'd2))}))});
  localparam [5:0] p8 = (~^(2'd0));
  localparam signed [3:0] p9 = {(4'd6),(3'sd1)};
  localparam signed [4:0] p10 = ((3'd4)?(5'd9):(2'd2));
  localparam signed [5:0] p11 = {(5'd27)};
  localparam [3:0] p12 = {(4'sd3),(-3'sd2),(5'd3)};
  localparam [4:0] p13 = (~|((((4'd2)^(4'd7))^~(&(2'sd1)))==={4{(5'd17)}}));
  localparam [5:0] p14 = ((5'd2 * ((2'd3)&&(4'd5)))||(((3'd5)?(4'sd0):(3'sd0))==(~^(-2'sd0))));
  localparam signed [3:0] p15 = (!(-(-5'sd9)));
  localparam signed [4:0] p16 = {(~|(!(2'sd0)))};
  localparam signed [5:0] p17 = (((+{(-2'sd0)})>=((5'd7)||(2'sd0)))===(4'd15));

  assign y0 = (~&(|(&{4{p3}})));
  assign y1 = (~^((a0-b2)?(~|a0):(p3?a5:b2)));
  assign y2 = (^((((&a2)<<(a3|b5))!={{a0,a0,p7}})<=(~&{(b5<=p11),(~(b3&a0))})));
  assign y3 = ((p12<<<p9)-(b1));
  assign y4 = (-(({p10,p17,b3}>>(p5!=p17))?({2{p1}}?{p0,p6,b0}:{p13,p14,p16}):{3{(p8?p7:p7)}}));
  assign y5 = (&({((-p4)?{p1,p1,p2}:(^p12)),$unsigned((~&(|(p16?p3:p15)))),({p4,p11}?(p8?p14:p11):{p10,p16})}));
  assign y6 = $unsigned(((4'sd6)===(5'd9)));
  assign y7 = ((a2?p13:b2)&&(p4?a2:b2));
  assign y8 = ((p10?b1:p12)?(^(b3?p5:b5)):(p14?p5:p16));
  assign y9 = {3{a5}};
  assign y10 = (^((2'd3)?{2{a0}}:(p5-a1)));
  assign y11 = ((((p13&&a0)==(a5|b1)))+(((a2>p15)<=(b4))||{(~p17),(!p0)}));
  assign y12 = ((&(4'd5))!=(4'd2 * (a0==a0)));
  assign y13 = (3'd3);
  assign y14 = (~^((~&(~|((b1^~b2)<=(b4?b5:a5))))<<({(a5-b2),(p10|a3)}<=((+b2)&&(a2?a0:a0)))));
  assign y15 = (~&({{a2,p2}}&&(p16>b0)));
  assign y16 = ($unsigned((~|(|$unsigned((~&(5'd2 * (p13*p0))))))));
  assign y17 = ((a3^p8)-(p6>>>p15));
endmodule
