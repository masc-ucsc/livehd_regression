module expression_00871(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(~|(((-5'sd7)>>>(3'd3))^{2{(2'd3)}}))}};
  localparam [4:0] p1 = {1{({4{(4'sd0)}}&&({3{(-5'sd1)}}-((3'd5)<<(4'd3))))}};
  localparam [5:0] p2 = (4'd1);
  localparam signed [3:0] p3 = ({4{(4'd4)}}?{1{{4{(4'd4)}}}}:{3{(3'd0)}});
  localparam signed [4:0] p4 = (6'd2 * (~|((5'd18)|(5'd25))));
  localparam signed [5:0] p5 = (+(5'd29));
  localparam [3:0] p6 = (-2'sd0);
  localparam [4:0] p7 = (+((4'd3)>=(3'd7)));
  localparam [5:0] p8 = (((4'd7)==(5'd29))&(~^(3'd0)));
  localparam signed [3:0] p9 = (((-2'sd0)&&(4'sd2))>>>(-4'sd5));
  localparam signed [4:0] p10 = {((((5'd19)>>>(-3'sd1))==={(4'sd3),(5'd0)})||((5'd10)!=(-(3'sd2)))),(~^((~{4{(-4'sd3)}})==((3'd1)>>>(5'sd11))))};
  localparam signed [5:0] p11 = (((5'sd6)?(5'd0):(5'sd4))&((3'd1)?(5'd7):(2'd2)));
  localparam [3:0] p12 = (2'd3);
  localparam [4:0] p13 = (-(&(~(&(~(-(&(~|(~&(~|(+(~(~&(5'd0))))))))))))));
  localparam [5:0] p14 = (~((4'sd2)<<<(-2'sd1)));
  localparam signed [3:0] p15 = {1{{4{((3'sd2)<(5'd28))}}}};
  localparam signed [4:0] p16 = ((4'd4)?{(~|(-4'sd7)),((3'sd2)<(-3'sd3))}:(3'd1));
  localparam signed [5:0] p17 = (~&(&((((-4'sd4)==(-4'sd3))>((2'd2)===(-2'sd0)))^~((+(5'd12))<<<(^(2'd1))))));

  assign y0 = ({(($signed((|{1{(~|$unsigned((a2<<p8)))}})))|{4{$unsigned(a1)}})});
  assign y1 = {({(a2==b5),(a2?a3:b5),(p11|a4)}|((p12?a5:a5)<<<(4'd2)))};
  assign y2 = {1{p5}};
  assign y3 = $unsigned((((3'sd3)>$signed(p14))?$unsigned((!(a2>=a4))):((b2+p12)?{2{p13}}:(5'd14))));
  assign y4 = {1{({{p4,p15,p3},{2{p6}}}-{{3{p5}},(p4&&p17),(p16|p13)})}};
  assign y5 = (($unsigned((p13?p9:p4))|((p15)+(p7?p5:p0)))<<<($signed($signed(p10))?(p6?p3:p4):(p5?p6:p1)));
  assign y6 = (((3'd4)?((p6>>>p10)?(p13?p0:p9):$unsigned(p4)):((6'd2 * p8)?(p10<<<p14):(2'd3))));
  assign y7 = {{4{{1{((a2?a3:b4)===$signed(b1))}}}}};
  assign y8 = (($signed($signed(p5))&&$signed($unsigned(p17)))>>>($signed((-b1))>>>(p2<<p12)));
  assign y9 = {(!(~|{a2,b4,p6}))};
  assign y10 = (p8^~p12);
  assign y11 = ({(-2'sd0),{4{a3}}}&&$unsigned($signed(($signed(($unsigned((4'd2 * a2))||(a2>=b5)))))));
  assign y12 = {((a4^~a0)<<<(6'd2 * a1)),((~&p17)>>(~|p9)),{{a2,a0,b1},(a5>>>b4)}};
  assign y13 = ((p11/p7)!=(p2%b1));
  assign y14 = (~|($unsigned((~^$unsigned((3'sd0))))));
  assign y15 = {(((^b4)+{3{a1}})&({a3,a4}&(a5===b4))),(({3{p4}}||(a3<<<a0))<={b1,a1,b2})};
  assign y16 = (a4==a2);
  assign y17 = ((({3{p1}}^~(~^p17))^((p12||p10)^~(~|p5)))<(^((p2>p9)==(p5!=p16))));
endmodule
