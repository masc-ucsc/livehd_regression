module expression_00684(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd1)*(5'd22));
  localparam [4:0] p1 = {4{{2{(-2'sd1)}}}};
  localparam [5:0] p2 = ((~^(~|(3'd1)))<<((3'd5)<=(4'd2)));
  localparam signed [3:0] p3 = (&(((3'sd0)?(2'd0):(3'd4))?((5'd13)?(5'sd11):(5'd12)):(~^{(2'd3),(2'd0)})));
  localparam signed [4:0] p4 = (~^(-(((+(2'sd0))>>>{(-2'sd1),(5'sd6)})?{(!(5'd8)),{3{(-4'sd1)}}}:(((4'd7)?(3'sd0):(-5'sd8))!=((2'd1)?(4'd15):(4'd12))))));
  localparam signed [5:0] p5 = ((5'sd5)<<<(4'sd5));
  localparam [3:0] p6 = (((2'sd1)+(-2'sd1))&&((-5'sd3)>(-5'sd4)));
  localparam [4:0] p7 = (((|(-4'sd5))?((-2'sd1)>>>(3'd4)):((2'd1)>=(4'd4)))===(((5'd12)>=(2'd2))?((4'sd1)==(5'sd10)):((4'd1)>>>(-5'sd10))));
  localparam [5:0] p8 = ((((-3'sd0)==(2'd2))>(3'd6))^(-((~^((2'd3)===(4'd0)))-(~^(~(5'd11))))));
  localparam signed [3:0] p9 = (!(!(-(-(^(3'd3))))));
  localparam signed [4:0] p10 = {{(2'sd1)},(-4'sd2),(5'd28)};
  localparam signed [5:0] p11 = (((5'sd12)?(3'd4):(3'd7))?{4{(3'd7)}}:(|{1{(4'sd2)}}));
  localparam [3:0] p12 = ((-3'sd3)<((5'sd1)==(5'sd9)));
  localparam [4:0] p13 = {3{(-(-{(-3'sd3),(5'd1),(-3'sd3)}))}};
  localparam [5:0] p14 = (&{{((3'sd0)^(-2'sd1))},(~|{(3'd4),(-3'sd0),(-4'sd7)})});
  localparam signed [3:0] p15 = (5'd3);
  localparam signed [4:0] p16 = (({(3'sd0),(3'sd3),(5'sd4)}?(~(2'sd0)):(~(4'd3)))?(~&((2'd2)?(3'sd1):(3'd5))):(~(5'd8)));
  localparam signed [5:0] p17 = {2{(5'sd10)}};

  assign y0 = {(~^(({(-{p15})}<<<((p16<<<b0)>(&p1)))&&(((-p7)|{a1,p8})^~{(p3<<b4),(b2>>>a1)})))};
  assign y1 = {3{{4{a1}}}};
  assign y2 = (~|{(5'd8)});
  assign y3 = {3{b0}};
  assign y4 = ((p15^b5)<<<(p1^p15));
  assign y5 = ({$signed(a0),(p1^p15)}>(5'sd11));
  assign y6 = ((a2>=b1)=={2{a0}});
  assign y7 = ({3{a3}}&{1{a3}});
  assign y8 = ({4{p0}}-({2{b1}}^~{3{p17}}));
  assign y9 = (~^(~&(((~a1))&&((a3||a3)))));
  assign y10 = (((a5===a4)?{1{(p10<<p11)}}:{1{(a0<=p11)}})-(((5'd2 * b1)!==(b2?b0:a3))-((a3>>b0)!=={3{a2}})));
  assign y11 = (6'd2 * (3'd6));
  assign y12 = ($signed((+$signed((p0?a2:p15))))!=(~|($signed((p10|p13))%p3)));
  assign y13 = {4{b4}};
  assign y14 = (^(3'd5));
  assign y15 = ($unsigned((a5?p14:p15))?$unsigned((&(b4>>>p6))):((b1?p11:a2)?(b0?p5:p11):(b5)));
  assign y16 = ((p11?p11:p8)?($unsigned(a3)<=$unsigned(b0)):{b0,b3,a3});
  assign y17 = ((-b2)?(a0?p13:b2):(&b1));
endmodule
