module expression_00645(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd5)&&(5'd5));
  localparam [4:0] p1 = ((-4'sd1)?(-3'sd1):(2'sd1));
  localparam [5:0] p2 = {4{(5'd15)}};
  localparam signed [3:0] p3 = (((3'd1)&(4'd0))&&((4'sd7)==(5'd15)));
  localparam signed [4:0] p4 = (!(2'd0));
  localparam signed [5:0] p5 = ({(~&{(-4'sd2),(3'd4)}),{{1{(3'sd2)}}}}+{1{{2{((-2'sd0)>(4'd14))}}}});
  localparam [3:0] p6 = (~((~&((~(4'd8))<=((5'd21)>(4'sd0))))>=((-3'sd1)+{(2'd1),(2'sd0),(3'd1)})));
  localparam [4:0] p7 = ((3'd0)%(-4'sd2));
  localparam [5:0] p8 = (((2'd3)>>>(4'd15))|{(-5'sd0)});
  localparam signed [3:0] p9 = {(~(-5'sd9)),(~&{1{{{(4'd12)}}}}),(5'd2 * ((3'd7)>(4'd1)))};
  localparam signed [4:0] p10 = {3{(((5'd9)^(2'd0))<<<((-3'sd3)?(5'sd0):(-3'sd1)))}};
  localparam signed [5:0] p11 = (~(4'd11));
  localparam [3:0] p12 = {(((-2'sd1)?(4'd13):(5'd26))?{2{(5'd2)}}:{4{(-3'sd1)}}),({(5'sd8),(-4'sd3)}<<<{4{(4'd15)}})};
  localparam [4:0] p13 = (((5'd24)<(2'd1))&&{(4'd15),(5'd31),(3'sd3)});
  localparam [5:0] p14 = (((^((5'd25)|(4'd12)))<=(^(~^(5'd8))))<=((~|((2'sd1)!=(4'd15)))<(!((3'sd0)<(-5'sd15)))));
  localparam signed [3:0] p15 = (|((5'd0)!==(4'd12)));
  localparam signed [4:0] p16 = ((~&{1{(!(4'sd4))}})&(|(!((3'sd0)!==(3'sd3)))));
  localparam signed [5:0] p17 = (((5'sd2)?((5'd15)*(-4'sd6)):(2'd1))^~(5'd17));

  assign y0 = ((+(|$signed($unsigned((a1!==b0)))))?($unsigned((p9%p9))==$unsigned((b2?a1:b1))):(((~|a2))==(4'd2 * p6)));
  assign y1 = $signed((5'd5));
  assign y2 = (~&((((p13?p16:a3)==(b0?p13:p1))>>(a2?p6:p6))<<<(~&(~&{{(p16?p11:p9)},(^(~&p1))}))));
  assign y3 = {(-4'sd5),(a0^~p7)};
  assign y4 = ((a1+b1)==(b2<<<a0));
  assign y5 = (((+(2'd2))||(-3'sd0))^(-3'sd3));
  assign y6 = (5'd2 * (+(|a2)));
  assign y7 = (((&$signed((p9+p0)))-((~b4)^~(~|p15)))>=((+(4'd2 * (p7-a0)))));
  assign y8 = (^(-4'sd3));
  assign y9 = (~|p15);
  assign y10 = (~((5'sd8)<=((4'sd5)&(3'd4))));
  assign y11 = ((-{3{b1}})?(|(a1?a3:a4)):$signed({3{a0}}));
  assign y12 = (((~^(6'd2 * b0))?(~|(a4&&a3)):(b5&&b5))===(-((^(a3&b0))<<<(~(b4?b3:b2)))));
  assign y13 = (~(&((4'd2 * (b2==b1))!=((b0-a2)!=(a1|b3)))));
  assign y14 = {(a1?b5:p14),(-3'sd0),(-5'sd2)};
  assign y15 = (((b2^~p9)-(p11&&p1))|((p9&p4)?{p2}:(p17>p9)));
  assign y16 = (5'd8);
  assign y17 = $unsigned((p3?a4:b0));
endmodule
