module expression_00576(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd3),(2'sd1),(3'sd2)};
  localparam [4:0] p1 = ((^(4'd2 * ((5'd13)<=(5'd0))))?{1{({2{(2'sd0)}}!=((-3'sd3)>=(3'sd2)))}}:(((-3'sd0)&&(3'sd1))<<<((2'd1)?(2'd2):(5'd2))));
  localparam [5:0] p2 = {2{({1{(~(4'd5))}}<<<((-4'sd2)>(3'd7)))}};
  localparam signed [3:0] p3 = (2'sd1);
  localparam signed [4:0] p4 = ({3{(~&(4'd1))}}^(~{1{(-2'sd1)}}));
  localparam signed [5:0] p5 = {{{(-3'sd3),(5'sd10),(4'sd5)},{(3'sd2),(5'd13),(3'd0)}},{{(2'd3),(3'd2)},{(-3'sd3)}},{{{{(4'd0),(4'd0)}}}}};
  localparam [3:0] p6 = ((-4'sd1)<(-3'sd2));
  localparam [4:0] p7 = (5'sd3);
  localparam [5:0] p8 = (4'd3);
  localparam signed [3:0] p9 = (((-4'sd7)>>(2'd0))+(3'd7));
  localparam signed [4:0] p10 = (5'd13);
  localparam signed [5:0] p11 = {{3{(4'd11)}}};
  localparam [3:0] p12 = ({(((2'd2)?(-4'sd4):(5'sd10))!=((3'sd1)?(5'd15):(3'sd2)))}>>>{((4'd7)?(4'd1):(3'sd3)),((3'd0)>>(2'd0))});
  localparam [4:0] p13 = ((-3'sd3)&&(^(3'sd0)));
  localparam [5:0] p14 = ((-5'sd4)?(5'd2 * ((3'd0)<<(4'd1))):(((-4'sd6)>>>(2'sd0))<<(-3'sd0)));
  localparam signed [3:0] p15 = (-(|(2'd3)));
  localparam signed [4:0] p16 = (~&(2'd0));
  localparam signed [5:0] p17 = (+((-((3'd5)^(5'sd4)))>(~|(!(4'd10)))));

  assign y0 = (3'd3);
  assign y1 = (&{2{({3{p11}}?(~^p17):(p2?a1:p13))}});
  assign y2 = ((p8&p10)<<{2{b3}});
  assign y3 = $unsigned((((^p10)*(~|p0))^~($unsigned(b1)!=(b5))));
  assign y4 = (p6?a0:a4);
  assign y5 = (~|((~(~|(a0?b5:b5)))?{4{p9}}:(((p13<<a3)))));
  assign y6 = (-3'sd3);
  assign y7 = ((p11+p15)<=(b5===b4));
  assign y8 = (((5'd13)<<{{b1},(~&p9)})+((5'd4)===((b0&b0)>>>(-4'sd4))));
  assign y9 = $signed(((((4'd2 * p14)?(p1?b1:a1):(b2|p12))?((a3||p17)?(a4?p3:b1):(p5*b4)):(~&((a0===a5)?(p3?p8:a5):(-p13))))));
  assign y10 = ((~((4'd13)?(p9|p7):(b0%p3)))<=((p5>a4)?(a2?b2:a1):(~b4)));
  assign y11 = (-(3'd7));
  assign y12 = ((b3?b1:a5)?(b3?a1:b4):(p9?a4:b1));
  assign y13 = {1{{2{(({4{p4}}&(4'sd0)))}}}};
  assign y14 = {a2,a5,p9};
  assign y15 = {$signed({1{(~|{2{(~|$unsigned((a0?a5:b1)))}})}})};
  assign y16 = ($signed((((p11<<b4)!=(a1*p5))>>>((a4-p12)||(a2==p12)))));
  assign y17 = (((b3?b4:a1)%b0)<<(~&(~((~&(a3?b5:b2))?(~&(^p1)):(b1&&a3)))));
endmodule
