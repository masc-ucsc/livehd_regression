module expression_00492(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{((!(2'd3))^~(~^(-4'sd7)))}}&&({((-4'sd6)&&(-5'sd14))}^~(~|{(-4'sd4),(3'd2),(3'sd2)})));
  localparam [4:0] p1 = (6'd2 * ((5'd20)!==(4'd14)));
  localparam [5:0] p2 = (5'd2 * (2'd3));
  localparam signed [3:0] p3 = {1{(-{4{(~{3{(-2'sd0)}})}})}};
  localparam signed [4:0] p4 = (2'd3);
  localparam signed [5:0] p5 = ((-(~((2'd3)&(2'd2))))||(~((-5'sd6)===(4'd14))));
  localparam [3:0] p6 = ({2{{(3'd0),(-4'sd5),(4'sd2)}}}<={(~^(5'd29)),((-5'sd7)?(5'sd12):(4'sd4)),((2'd0)>>>(3'd4))});
  localparam [4:0] p7 = ((5'd18)<=(2'd3));
  localparam [5:0] p8 = ((((3'sd3)&(3'sd3))<<((5'sd13)===(3'sd0)))||(~^(|(((4'd14)>(2'd2))>>>((2'sd1)||(3'd1))))));
  localparam signed [3:0] p9 = (5'd3);
  localparam signed [4:0] p10 = ((2'sd0)+(2'd0));
  localparam signed [5:0] p11 = ((((3'sd3)?(3'd6):(5'sd8))<((~^(3'sd3))^~((2'd3)===(5'd23))))|{4{{2{(3'd5)}}}});
  localparam [3:0] p12 = (((((2'd2)&&(-4'sd3))||(^(2'sd1)))|((~&(2'd3))+((2'd1)==(2'd2))))===(!(((4'sd6)+(4'd2))<<((2'sd0)<(2'sd1)))));
  localparam [4:0] p13 = (((4'd6)?(3'd5):(-5'sd1))<=(!((-4'sd0)==(3'd5))));
  localparam [5:0] p14 = {1{{(5'sd2),(5'd19)}}};
  localparam signed [3:0] p15 = (4'd10);
  localparam signed [4:0] p16 = (~&({4{((3'sd2)<(2'd0))}}&&(~(~{2{(~^(4'd3))}}))));
  localparam signed [5:0] p17 = ({{(-4'sd3),(4'd5),(3'd7)}}>>>{(-2'sd0),(5'd0),(5'sd9)});

  assign y0 = (~^{2{{3{b4}}}});
  assign y1 = (5'sd9);
  assign y2 = {((b4?b4:b2)==={a3,b3,a0}),((b0>a5)?(a0?b0:p1):(^p5)),((b5?b0:p0)||(p8<p4))};
  assign y3 = (~^{b4});
  assign y4 = (|((p12?b2:p2)?(-(~p9)):(p7?b1:p4)));
  assign y5 = {$unsigned(((-4'sd7))),(4'd7)};
  assign y6 = (!(-2'sd0));
  assign y7 = {(!({(p0-p5),(5'd2 * p0),(p11>>p0)}>=(-5'sd6)))};
  assign y8 = (((~|p5)?{p15}:(p11?p0:a3))?{{p9},(p10),$signed(b1)}:(~^(~(~(&p10)))));
  assign y9 = (6'd2 * {b0,p2,a0});
  assign y10 = (({(a0^a0)}?(a1|a1):(b4<b5))===(3'sd0));
  assign y11 = (((&(p1?p2:p0))<<<((p13^~p6)?(p5?a5:p15):(p8?p10:p6)))==(5'sd13));
  assign y12 = ((|p4)?(6'd2 * p13):(b4===a0));
  assign y13 = (3'd4);
  assign y14 = {3{{{a5},{3{b0}}}}};
  assign y15 = (5'd4);
  assign y16 = (3'sd3);
  assign y17 = (~^($unsigned(((p7-p0)/a3))?((a2^a2)===$signed((a4))):(3'd2)));
endmodule
