module expression_00738(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd0)&(~|(~^((+(3'd1))<<(~(3'd6))))));
  localparam [4:0] p1 = (2'd2);
  localparam [5:0] p2 = (6'd2 * ((4'd5)>=(5'd4)));
  localparam signed [3:0] p3 = {4{{3{(-3'sd1)}}}};
  localparam signed [4:0] p4 = {3{(3'd3)}};
  localparam signed [5:0] p5 = {(4'd12),(3'd3)};
  localparam [3:0] p6 = ((((4'd13)<(-2'sd0))^~{(-5'sd10),(5'd2),(-3'sd1)})?{(2'd3),(2'd2),{(4'd10),(3'sd3)}}:((5'd29)?(2'd2):((4'sd5)?(-4'sd6):(-3'sd0))));
  localparam [4:0] p7 = ((4'd13)>(4'sd1));
  localparam [5:0] p8 = {4{(~|(-4'sd5))}};
  localparam signed [3:0] p9 = {((&((5'd8)&(5'd17)))>=(((3'd6)?(5'd9):(5'd30))!=={(-2'sd1),(-3'sd2),(4'd12)}))};
  localparam signed [4:0] p10 = ((((3'd6)<<(4'sd0))^~(~(4'sd7)))<<(((-5'sd15)|(3'd7))+((-4'sd6)>=(4'd7))));
  localparam signed [5:0] p11 = (|((3'd0)-(3'd5)));
  localparam [3:0] p12 = (3'd4);
  localparam [4:0] p13 = (~|(+(^((|(3'd5))||((5'd17)>>(-4'sd0))))));
  localparam [5:0] p14 = (((3'd6)+(3'd4))^~((2'd1)^~(-2'sd0)));
  localparam signed [3:0] p15 = ((((5'd23)&&(4'd5))>=((2'sd0)^(3'd2)))<<<(!(&((5'd23)^~(4'sd6)))));
  localparam signed [4:0] p16 = (|((5'sd10)&&(4'sd1)));
  localparam signed [5:0] p17 = {4{(-2'sd1)}};

  assign y0 = (~({4{{4{b2}}}}>>>((p16>>p10)==(+(~^b1)))));
  assign y1 = ((4'd1));
  assign y2 = ((a3!==a4)<<<(b1^a5));
  assign y3 = ((~&(|(5'sd14)))<((5'd14)|(~|(4'd7))));
  assign y4 = ({4{(p1<=p6)}}==({(b3<<<a2),(~&p5)}>>(+{3{p0}})));
  assign y5 = {p3,p5};
  assign y6 = {3{{{p10,b5,p0},{4{b2}}}}};
  assign y7 = ((4'd2)|(-2'sd0));
  assign y8 = {1{($signed((4'd3))^~{3{(p2&p17)}})}};
  assign y9 = {2{(2'd2)}};
  assign y10 = ({{p3,p12,b3},(b5==a4),(~|(a3?p14:b0))}==({(~^{b2,a0})}^~(b5?p17:b0)));
  assign y11 = (({(a2^a2)}<<<{(p17>>>b4)})>=(({a2,a1}<=(b0<a4))||((a0!==b4)+(b0>>b2))));
  assign y12 = (-(~|((((^b2)!=(b5>>>a1))^~((a5>>>a0)&&(^a3)))===(~|(~|(-(+((~&a5)<(^a4)))))))));
  assign y13 = (((~(+b1))===(b3^b4))<=(^((-b5)!=(a1-b3))));
  assign y14 = (|a1);
  assign y15 = $signed({4{(b5^~b0)}});
  assign y16 = ({1{(~|(!{2{(-a2)}}))}}>>>((&(~&p17))&(^(a3^~a0))));
  assign y17 = (&(+(((a1^~a2)+(&p12))>>>((b2?a5:p8)||(p14?b4:b2)))));
endmodule
