module expression_00379(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{(-2'sd1)}}+(~|(2'sd0)));
  localparam [4:0] p1 = {1{(2'd0)}};
  localparam [5:0] p2 = (^{1{(3'd5)}});
  localparam signed [3:0] p3 = {3{(((5'd7)===(3'd5))|((-5'sd3)?(2'sd0):(5'sd6)))}};
  localparam signed [4:0] p4 = ({1{(|(((-4'sd5)<<(5'd12))&{3{(-2'sd1)}}))}}+{2{({3{(4'sd4)}}||((-5'sd6)>>>(5'd19)))}});
  localparam signed [5:0] p5 = {(4'd12),(4'd2),{(-5'sd1),(-4'sd1)}};
  localparam [3:0] p6 = ((2'd3)<=(((3'd3)||(3'd6))%(5'd14)));
  localparam [4:0] p7 = ((((5'sd3)>>>(-2'sd1))*((5'sd1)?(5'sd3):(5'sd13)))<=(((3'd2)?(4'sd4):(-4'sd7))?((-5'sd13)>>>(4'd10)):((3'sd1)^~(3'd2))));
  localparam [5:0] p8 = {(-5'sd15),((+(3'd6))<(^(4'sd2))),(((4'sd1)?(3'sd3):(-4'sd4))&&(~^(5'd5)))};
  localparam signed [3:0] p9 = (((&((2'd2)%(4'd11)))>=((4'sd1)!==(3'd7)))|((&((4'd15)===(3'sd0)))||((4'd2)<(-3'sd3))));
  localparam signed [4:0] p10 = (((-2'sd1)/(4'sd4))?(6'd2 * (3'd5)):((2'sd1)<=(-5'sd12)));
  localparam signed [5:0] p11 = (-(~&(~&(-((-(2'sd1))?(^(5'd31)):(~^(4'sd2)))))));
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = (~(2'sd1));
  localparam [5:0] p14 = ((-4'sd3)^~(2'sd0));
  localparam signed [3:0] p15 = (^((5'd4)>>(+(5'sd7))));
  localparam signed [4:0] p16 = {{1{{(4'sd7)}}},{(3'sd3),(-4'sd6),(3'd0)},{1{{2{(3'sd0)}}}}};
  localparam signed [5:0] p17 = {{{{((4'd3)?(4'd3):(4'd1))}},{(!(5'd9)),(^(4'd5))}}};

  assign y0 = (~|{2{{1{a2}}}});
  assign y1 = (4'd2);
  assign y2 = (4'd14);
  assign y3 = (~((~&b0)&(b2!=p2)));
  assign y4 = (((p3==p8)^~(p16?p1:p4))<={3{(p12^~p11)}});
  assign y5 = ($signed((-2'sd1))>>>((^(-(b2||p6)))&$signed((a2<p15))));
  assign y6 = $signed($unsigned((((p14/b5))%p17)));
  assign y7 = {1{(~&({2{p9}}>{3{p11}}))}};
  assign y8 = ((|((|(p8?a0:a5))?(|(-p14)):(b2>p13)))!=(~^(+((+(~^(!p13)))<(~|(!(|p2)))))));
  assign y9 = ({(p2>=b1),(p1),(b4<<b4)}>>$signed(((p12-b2)<<<$unsigned(b5))));
  assign y10 = (((b5>>>p1)<(p7?p7:b0))&&((p13>p3)==(p11+p4)));
  assign y11 = ((-5'sd1)?(p9?p3:b4):(4'd2));
  assign y12 = (((p9?a5:p16)==(2'd0))&(((5'sd5))!==(-5'sd5)));
  assign y13 = $unsigned((4'd6));
  assign y14 = (((p10^a1)>>(p17>>>a5))^~(5'd2 * (a1!==b0)));
  assign y15 = {2{((+b3)?{1{p0}}:(4'd2 * b1))}};
  assign y16 = (-((b0>>>b2)|(4'd2)));
  assign y17 = ((((b2)&&(3'sd0))&&({2{b4}}-(b3!=p6))));
endmodule
