module expression_00135(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-4'sd7)|(-2'sd0))<<<((2'sd1)+(4'd11)));
  localparam [4:0] p1 = (((-2'sd1)!==(-2'sd1))==(5'sd11));
  localparam [5:0] p2 = (~((!(5'd8))==(~|(4'd10))));
  localparam signed [3:0] p3 = (((+(~^(3'd2)))==(~((2'd2)!=(5'd11))))===((~&((5'd7)^~(5'd11)))<=(^(~&(4'd8)))));
  localparam signed [4:0] p4 = (2'sd1);
  localparam signed [5:0] p5 = ((-3'sd0)?((2'd0)?(5'sd5):(-3'sd0)):{4{(4'd14)}});
  localparam [3:0] p6 = ({(4'd0),(3'sd3),(-4'sd3)}?(~^(-3'sd2)):(^(3'd6)));
  localparam [4:0] p7 = (-3'sd2);
  localparam [5:0] p8 = ((3'd1)<<<((5'sd15)?((3'sd3)?(4'd15):(-2'sd1)):((-2'sd1)&&(3'sd3))));
  localparam signed [3:0] p9 = ((5'd2 * (5'd28))=={3{(-2'sd0)}});
  localparam signed [4:0] p10 = (4'sd4);
  localparam signed [5:0] p11 = ({(~|(-3'sd1)),((-4'sd0)>=(-3'sd2)),(|(3'd1))}<(~^({(-5'sd0),(5'd0),(-3'sd2)}>(+(3'd2)))));
  localparam [3:0] p12 = (3'd3);
  localparam [4:0] p13 = {(2'sd1)};
  localparam [5:0] p14 = (((4'd7)/(3'd6))>(2'd0));
  localparam signed [3:0] p15 = (+((2'd1)^(2'sd1)));
  localparam signed [4:0] p16 = {(|{(~(5'sd5)),{(5'sd11),(3'd2),(3'd2)},(-(4'sd7))})};
  localparam signed [5:0] p17 = ((2'd3)^(-4'sd6));

  assign y0 = $signed(({1{{1{((p4|p17)!=(p16?p3:p15))}}}}!={4{(4'd2 * p8)}}));
  assign y1 = {p6,p11};
  assign y2 = {1{(p15>=p10)}};
  assign y3 = (-$unsigned((!{1{$unsigned(({3{(~&a1)}}&$unsigned((~|{4{b5}}))))}})));
  assign y4 = (+(5'sd5));
  assign y5 = (~&((|(({1{a5}})^~{2{b1}}))<<<(~(~&({2{p9}}+(b0<a3))))));
  assign y6 = {1{($unsigned(((p6>>>p15)>>(p9!=a1)))=={3{$unsigned(p12)}})}};
  assign y7 = {4{{4{p0}}}};
  assign y8 = $unsigned((-((4'd3)+(p6==p9))));
  assign y9 = (!{4{$unsigned(p1)}});
  assign y10 = $signed((-5'sd11));
  assign y11 = (!(-4'sd0));
  assign y12 = (|{({p10,p6,p8}&&(p12==p12))});
  assign y13 = {3{(a1?p8:a4)}};
  assign y14 = ({4{{3{b0}}}}?{3{(p13<<<p9)}}:((p3?p15:p6)?(5'd2 * b1):(p10?p13:p12)));
  assign y15 = ($signed(((4'sd0)>>>(-3'sd2)))?((b0!=p8)<(p11||p4)):(&{(2'sd1)}));
  assign y16 = {4{(&(p16&a3))}};
  assign y17 = (&{(^(^(~|{{a2},{b3,a0}}))),{{(|{(~&a2),{p17,a1},{p1,p17}})}}});
endmodule
