module expression_00365(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'd3)^(4'd0))!=((3'd1)===(-3'sd1)))>>(((3'd1)<(-5'sd0))-(~&((4'd0)^~(-5'sd14)))));
  localparam [4:0] p1 = ((4'sd7)&&(-2'sd0));
  localparam [5:0] p2 = {1{((|(~^{2{((4'sd4)^(5'sd5))}}))!=({2{(2'd2)}}-(6'd2 * (3'd7))))}};
  localparam signed [3:0] p3 = (((5'd15)?(3'd6):(2'd2))?((5'd23)&&(2'sd1)):((-2'sd0)%(3'd2)));
  localparam signed [4:0] p4 = (-(!(~^(~&(&(~^(-(|(+(~|(~(~(-2'sd1)))))))))))));
  localparam signed [5:0] p5 = ({(-2'sd1),(2'd0),(-3'sd1)}?(3'd2):(!{(-4'sd2),(4'd2),(5'sd10)}));
  localparam [3:0] p6 = (((4'd11)?(2'd2):(-4'sd2))-((2'sd1)>>>(3'd3)));
  localparam [4:0] p7 = (-2'sd1);
  localparam [5:0] p8 = (((3'sd0)>=(5'sd1))?((2'sd0)^(5'd30)):(2'd2));
  localparam signed [3:0] p9 = ((2'sd1)<<(5'd11));
  localparam signed [4:0] p10 = ((!(2'd0))?(4'd2):({(3'd0),(3'd2),(3'sd2)}<<(2'sd1)));
  localparam signed [5:0] p11 = (-((5'd16)<=(-(-3'sd3))));
  localparam [3:0] p12 = ((!((5'd29)?(-4'sd6):(5'sd0)))>>(~|((5'sd3)^~(5'd25))));
  localparam [4:0] p13 = ((((3'd0)<<<(2'd0))!=(-2'sd1))>>>(-5'sd3));
  localparam [5:0] p14 = ({3{((-5'sd4)>=(4'd15))}}!==((^(4'd0))>>((-5'sd5)?(2'd3):(4'sd6))));
  localparam signed [3:0] p15 = (|(4'd3));
  localparam signed [4:0] p16 = (5'd17);
  localparam signed [5:0] p17 = ({4{(-4'sd4)}}<((5'd7)<(2'd2)));

  assign y0 = ((((5'd31)&&(5'sd1))-((a3-a0)===(b5>>a3)))>>(2'd3));
  assign y1 = {((~|p3)?(&a5):(!p2))};
  assign y2 = (|(5'd2 * (a0?b0:a0)));
  assign y3 = (&(3'd2));
  assign y4 = ((p4?p8:p11));
  assign y5 = ((b0!=a0)*(b4*a0));
  assign y6 = {(((!b1))?(^(~p15)):{{a3}})};
  assign y7 = ({b5,p2,b4}<<<{(p15^p17)});
  assign y8 = (p13%p7);
  assign y9 = ((|((b5?a1:a1)<<<($unsigned(a4)>=(a3>>b2))))!==(((b2|a4)&&(b5===b0))==={4{a0}}));
  assign y10 = (((a4?b3:a2)?$unsigned(a0):(b1?b5:a0))?((a2?a4:b5)?(p13?b5:a3):(b1)):$unsigned((b0?p2:b1)));
  assign y11 = ($signed((((p10^a4)?$signed(p11):(a3<<<a5))))>(~^((p13>>b5)?(p7?p17:p8):(p4&b5))));
  assign y12 = ((6'd2 * (b2&&a2))>(3'd7));
  assign y13 = ((~^({1{$signed(b3)}}>>(-$signed(b4))))-(($unsigned(a4)&{4{a4}})>>>($unsigned(b3)^(p1<<<a5))));
  assign y14 = {(-5'sd9),$signed(p11),(4'd15)};
  assign y15 = (({{p17,p1,p6},(a4>>p5),((4'd2 * p6))})!={($unsigned({b3,b4,a4})!==$unsigned($unsigned({b4,a3,b1})))});
  assign y16 = (~^{4{(^(~&{3{p15}}))}});
  assign y17 = (({3{a0}}-((b2<=b1)===(a1-a5)))&{({(b3>>a1)}),((~|(~^p1)))});
endmodule
