module expression_00735(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-5'sd7)<<(2'd0))>((3'd6)>>(4'd12)));
  localparam [4:0] p1 = (((-2'sd1)<<(2'sd1))>=(~^(+(-2'sd0))));
  localparam [5:0] p2 = {((5'sd14)|(-2'sd0))};
  localparam signed [3:0] p3 = (((5'd24)>((3'd6)||(2'sd1)))^{((3'd5)-(-2'sd1)),{(3'sd3),(3'd6),(5'd16)}});
  localparam signed [4:0] p4 = (~(-4'sd2));
  localparam signed [5:0] p5 = (((4'sd3)<<(4'd1))-{{2{(2'd0)}}});
  localparam [3:0] p6 = (((5'd9)+(4'd13))?(~|(-5'sd8)):((3'd0)>=(-3'sd2)));
  localparam [4:0] p7 = ((5'sd15)&(4'd11));
  localparam [5:0] p8 = ((4'd0)!==((-3'sd3)!=(5'd23)));
  localparam signed [3:0] p9 = {((^(4'sd5))<(4'd9)),(!(^(2'd0)))};
  localparam signed [4:0] p10 = ({(3'd6),(3'd5)}!=={(3'd7),(4'sd5),(3'd3)});
  localparam signed [5:0] p11 = (!({(-3'sd2),(-3'sd3)}&((3'd6)-(-2'sd0))));
  localparam [3:0] p12 = {3{(-2'sd0)}};
  localparam [4:0] p13 = (^{2{(&(-3'sd3))}});
  localparam [5:0] p14 = ((|(^(3'sd0)))^(&{(4'd15),(4'd5),(2'd1)}));
  localparam signed [3:0] p15 = (!((~&(~&((-2'sd0)?(4'd2):(4'd14))))?(-3'sd1):(~&(&(~(2'd2))))));
  localparam signed [4:0] p16 = (^(4'd12));
  localparam signed [5:0] p17 = ((((&(3'sd0))==((5'd11)?(4'd12):(4'd11)))>((5'd0)?(5'd29):(4'd4)))!==(~|(|(~(~&(!((-2'sd0)^~(3'sd2))))))));

  assign y0 = ((5'sd8)&&(5'd18));
  assign y1 = (3'sd3);
  assign y2 = ({1{(p2|a2)}}>{(-4'sd5),{1{p13}}});
  assign y3 = ((p3<p13)?(a3>>>p14):(5'sd10));
  assign y4 = {p11};
  assign y5 = {((p2?p1:p17)&&(p1&p10)),{{p11},(b4<<<p3),{4{a0}}},({b4,p8}?(a4?p12:b5):{2{p6}})};
  assign y6 = (((p2<a4))?(~|{2{b5}}):(^(p5^~a1)));
  assign y7 = ({(a3?b4:a4),(b2||b3)}<<{{{a2,b0,b5}},(!{a0,b3})});
  assign y8 = ((p13>=p0)?(5'd13):(5'd23));
  assign y9 = (|(4'd2));
  assign y10 = (((a3===b1)&&(a1!=b3))&&(5'd2 * (b2&a0)));
  assign y11 = (((p13/a3)-(p14>=p16))-($unsigned($unsigned(a0))<=(b5<=p2)));
  assign y12 = ((-4'sd2));
  assign y13 = $signed(((b0)==(p14||a4)));
  assign y14 = ($unsigned((b1>>>b2))-{a4,b0,b4});
  assign y15 = ((~|{$unsigned({{b3,a3,p7},(-3'sd2)})})^(~&(((p14<p0)<<(a4))-(!(a0!==b0)))));
  assign y16 = (!{2{{{(|p7)},(-(~&p4)),(^(^b1))}}});
  assign y17 = {(&($signed(p16))),((+b0)>=(b1>>a0)),((a3===b1)-{a5})};
endmodule
