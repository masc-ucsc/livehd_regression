module expression_00706(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{((5'd25)<<<(-2'sd1))}};
  localparam [4:0] p1 = (6'd2 * ((4'd2)>=(4'd3)));
  localparam [5:0] p2 = {(2'd3)};
  localparam signed [3:0] p3 = ({(2'd2),(4'd8),(5'sd9)}===((4'd14)<<(5'd9)));
  localparam signed [4:0] p4 = ((-3'sd2)?(3'd3):(-2'sd1));
  localparam signed [5:0] p5 = ((((3'd6)!=(-5'sd7))||(&(2'd1)))||{4{(-5'sd2)}});
  localparam [3:0] p6 = (4'd0);
  localparam [4:0] p7 = ({2{(3'd5)}}>=((-4'sd3)?(3'd7):(5'd25)));
  localparam [5:0] p8 = (((-2'sd1)<<<(2'sd1))|((3'd3)|(-3'sd1)));
  localparam signed [3:0] p9 = (({{(4'd8)}}>{{(2'd0),(-3'sd1)}})<<{(((5'd4)-(5'd20))&{(-5'sd7),(5'd9)})});
  localparam signed [4:0] p10 = (((-5'sd6)<=(4'sd2))&&(5'd28));
  localparam signed [5:0] p11 = (~|(^(~|{1{(-{1{(&(4'd7))}})}})));
  localparam [3:0] p12 = {(|{((-5'sd14)?(2'd1):(-5'sd8)),(|(~(2'sd0)))})};
  localparam [4:0] p13 = (~&(~&(((5'd13)?(-4'sd6):(5'd7))?((-3'sd2)?(2'd1):(2'd2)):(|((-4'sd3)?(3'd5):(-2'sd0))))));
  localparam [5:0] p14 = (!(~&({((3'sd2)|(2'sd1)),((5'd1)||(5'sd9)),{(3'sd0),(4'd11),(3'd4)}}+(^(3'd0)))));
  localparam signed [3:0] p15 = (5'd10);
  localparam signed [4:0] p16 = {(-4'sd7),(4'd12)};
  localparam signed [5:0] p17 = (!(+(~&((3'd5)?((-5'sd3)?(4'd5):(4'sd2)):(4'd0)))));

  assign y0 = (~(^(5'sd4)));
  assign y1 = (~|((4'd2 * (p12^p7))-((a0&p13)?(p2<<<a0):(b0==p15))));
  assign y2 = ((-3'sd3)!=(&(!(+((p1!=a2)||(a3>>a0))))));
  assign y3 = $unsigned(b2);
  assign y4 = ((-((p0<<p11)^~(^p9)))-((p9+p13)&(p12||p11)));
  assign y5 = {4{{2{{1{p7}}}}}};
  assign y6 = $signed($signed((($signed((p0?p3:p16))))));
  assign y7 = (-3'sd3);
  assign y8 = {(~^(p13!=b2))};
  assign y9 = {$signed({b5,a3,a3}),(!(+p3)),(^(4'd5))};
  assign y10 = {({(b4?b4:b0),(p8?a4:a4)}?((5'd18)<(p0?b0:b1)):((b3&a0)!==(b3>>>a3)))};
  assign y11 = ((({a0,a3}!=={b5})>=((6'd2 * p7)<<(p15<<<p9)))+{({p0}-(a4===b3)),{(p3^~p6),(p8>>p12),(p9+p7)}});
  assign y12 = {((|(a2^b0))&{a0,a2,p5})};
  assign y13 = (&(~|(3'd4)));
  assign y14 = (($unsigned($signed(p15))&&(&(p16?p10:a1)))|$signed(((+p17)^~(a1?p9:p11))));
  assign y15 = ((a4^p16)<<<(!a2));
  assign y16 = ((2'd0)?(-4'sd7):((p16?p3:b5)?{1{b4}}:(3'd7)));
  assign y17 = {3{((a3?b1:p5)<<(b4>b1))}};
endmodule
