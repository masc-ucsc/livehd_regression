module expression_00349(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'd2);
  localparam [4:0] p1 = (-(|{4{(6'd2 * (2'd1))}}));
  localparam [5:0] p2 = ({{(2'sd0),(3'd7),(-3'sd1)},{(2'd2),(2'sd0),(2'd1)}}^{{(&(4'sd2)),((4'd5)&(4'sd1))}});
  localparam signed [3:0] p3 = ((5'sd6)==(3'd1));
  localparam signed [4:0] p4 = {{((3'd7)==(-2'sd0)),((-3'sd0)?(4'd13):(4'sd6)),((-3'sd1)?(-3'sd3):(2'd3))},({(5'sd8),(5'd27)}?((3'd5)?(2'd0):(4'd13)):{(4'd14),(5'd13)}),(((2'd3)==(2'sd1))>>((5'd3)>>>(2'sd0)))};
  localparam signed [5:0] p5 = (((5'sd13)?(-3'sd3):(5'sd1))?(+((2'd3)%(4'd2))):((2'd1)?(-3'sd1):(3'd0)));
  localparam [3:0] p6 = ((~(^(2'sd0)))<=((4'sd4)+(-5'sd5)));
  localparam [4:0] p7 = (|{{(-2'sd0),(3'd0),(2'sd0)},((-3'sd1)<(-2'sd0)),((4'sd4)>>>(4'd15))});
  localparam [5:0] p8 = {(((4'd7)!=(4'd12))^~((2'd2)||(-2'sd0))),({(5'd6),(-3'sd0),(4'd2)}<{(5'd13),(3'sd2),(5'd7)}),({(3'd5),(4'sd0)}<<((-4'sd7)^~(5'd4)))};
  localparam signed [3:0] p9 = ((((4'd0)/(5'd29))%(4'd8))>=(6'd2 * ((2'd0)<<<(2'd1))));
  localparam signed [4:0] p10 = {1{(2'd2)}};
  localparam signed [5:0] p11 = ({(4'sd7),(2'd2)}?((4'sd0)-(2'd3)):((5'd0)?(-5'sd12):(4'd14)));
  localparam [3:0] p12 = (|(&(-((((-2'sd1)^~(3'd4))<(~&(~|(-2'sd1))))<<(-(~^(-(&(!(-2'sd1))))))))));
  localparam [4:0] p13 = {(5'd2 * ((5'd27)?(2'd1):(2'd2))),(3'd1)};
  localparam [5:0] p14 = (~^(3'd3));
  localparam signed [3:0] p15 = (({4{(5'd7)}}?{4{(5'd2)}}:(-4'sd3))?({4{(5'd13)}}?(5'd2):((-3'sd3)?(-3'sd3):(2'd1))):{4{(2'd1)}});
  localparam signed [4:0] p16 = ({(4'd14)}&((4'sd1)==(5'd27)));
  localparam signed [5:0] p17 = ({(-4'sd2)}?((4'sd1)<<<(3'sd0)):((4'd8)!==(5'd30)));

  assign y0 = ((p11?b1:b2)?(&(~|b2)):(p1?a3:a3));
  assign y1 = (((p16!=p13)<<<(|p15))<<<((~^b4)!==(a1^~b2)));
  assign y2 = {{{(!(2'd3))}}};
  assign y3 = (|(-5'sd3));
  assign y4 = ((-4'sd3)==={3{{2{b0}}}});
  assign y5 = (((b3^~a4)^~(a2<=a5))?(-(4'd1)):((b0>b5)!=$signed((-2'sd0))));
  assign y6 = (2'd3);
  assign y7 = (~(5'd2 * (~|{p6})));
  assign y8 = (4'sd7);
  assign y9 = ({p2}||{a4,p13});
  assign y10 = {({p6,a3,p8}>(p4==b1)),{(6'd2 * p1),{p0,p11},{p5,p12}},((6'd2 * p1)>>>(p12||p11))};
  assign y11 = (&{1{{((^{(+p10),(~^p12),{3{p8}}})>={3{(&p16)}})}}});
  assign y12 = ({(p4==p15)}?(p12?p13:a3):(-3'sd3));
  assign y13 = (4'd2 * (~{3{b0}}));
  assign y14 = ((^$unsigned((({(p10==a1)}>=$signed((&b1)))))));
  assign y15 = ($unsigned({3{{3{p1}}}}));
  assign y16 = ((~^((3'd2)))<(~|(|((+(a1^~p8))?$signed((p13<<<p2)):(~(b1!=a0))))));
  assign y17 = ($signed((b3^~b3))!==(^(a3>>b3)));
endmodule
