module expression_00604(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-3'sd2)>>>(3'd3));
  localparam [4:0] p1 = ((6'd2 * ((4'd9)?(5'd21):(4'd6)))<(4'd15));
  localparam [5:0] p2 = (|(!(-4'sd1)));
  localparam signed [3:0] p3 = {1{{((-2'sd0)!==(5'd17)),((-2'sd0)!==(4'd6)),{(2'sd1)}}}};
  localparam signed [4:0] p4 = (-{{(3'd5),(5'd15)},(~^(-3'sd2)),((5'sd5)?(2'd3):(3'sd2))});
  localparam signed [5:0] p5 = (-((-5'sd5)^(-4'sd3)));
  localparam [3:0] p6 = ((((4'sd3)===(5'sd12))||{(^(5'sd10))})===(~({(5'd8),(-4'sd7),(3'd1)}||{(-4'sd7),(2'd2),(3'd4)})));
  localparam [4:0] p7 = (!(-4'sd6));
  localparam [5:0] p8 = ({((3'sd2)?(-3'sd3):(-5'sd3))}&((2'd3)?(-4'sd2):(-5'sd11)));
  localparam signed [3:0] p9 = ({((5'd4)<<<(3'd0)),((-3'sd2)?(2'sd0):(3'd1)),{(-3'sd2),(-3'sd3),(5'd22)}}<<(|{(((5'd28)?(2'sd0):(-5'sd7))?{(5'd13)}:(5'd15))}));
  localparam signed [4:0] p10 = (+((~&((4'd12)?(4'd0):(4'sd0)))?((~(3'd4))?(+(4'd6)):((-5'sd11)?(5'd14):(-4'sd5))):(|(~&(~&((3'd2)?(5'd1):(3'd6)))))));
  localparam signed [5:0] p11 = (-4'sd3);
  localparam [3:0] p12 = ({2{(3'sd2)}}?((5'd27)?(4'd3):(5'd17)):((-3'sd3)>>>(-2'sd1)));
  localparam [4:0] p13 = ({1{(4'd7)}}>{4{(5'sd12)}});
  localparam [5:0] p14 = (((+(4'd10))^~(~(-4'sd4)))>=(~|(~&((-4'sd0)-(2'd1)))));
  localparam signed [3:0] p15 = (({(2'd2),(5'd5)}|{(3'sd2),(-5'sd15)})^~({((-4'sd0)&&(-4'sd5))}==((3'd7)?(4'd7):(5'd6))));
  localparam signed [4:0] p16 = (-{3{(~|(((2'sd1)<<<(5'sd1))<(^(2'd3))))}});
  localparam signed [5:0] p17 = (~&(&(^(5'sd14))));

  assign y0 = (((~&{4{p8}})|(p7>>p13))^(5'sd10));
  assign y1 = ({3{b1}}<(-2'sd1));
  assign y2 = ($unsigned(({b4,a5}?{b3,p10}:{a0,b4}))!={{a3,b0,a4},(p1?a5:a1),$unsigned({p9,a5})});
  assign y3 = {2{(p8?b3:p13)}};
  assign y4 = {((a1?p11:p0)<<(a4-p8)),((p14?b4:a0)?(b0?p10:p5):(b1<<<b2)),((b1|a0)>(p15^p17))};
  assign y5 = (~&(^$unsigned((b2-p17))));
  assign y6 = {2{(~p15)}};
  assign y7 = ((((a3^~b3)>>(b3-b5))<<<((a1^~p6)-(~&b4)))+{(4'd2 * (|p13)),{(!a3),(+b4)}});
  assign y8 = {1{(~&(~|(((a3+b5)||{3{b2}})|{(~&p7),$signed(p12),(~p8)})))}};
  assign y9 = ((a5?a3:p8)?((&b1)<={1{b4}}):{(~|{4{b2}})});
  assign y10 = {1{{3{({b4,b3}&$signed({a1,b1}))}}}};
  assign y11 = ((|(4'd14))-(|(!$signed((-({p6,a3}^(-5'sd11)))))));
  assign y12 = ((2'd0)<<<{1{((-3'sd3)&&{4{p8}})}});
  assign y13 = (5'd6);
  assign y14 = (-(!(5'd3)));
  assign y15 = {2{((~&(~b5))?{2{a4}}:{2{a5}})}};
  assign y16 = $unsigned((a4?a3:a5));
  assign y17 = ({($unsigned(a4)||{b2})}!==((a5)==(b5)));
endmodule
