module expression_00747(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~^(4'd2))?((-3'sd2)||(3'd3)):((4'd12)+(4'sd2)))<(((2'sd1)%(5'd2))|(4'd2 * (3'd4))));
  localparam [4:0] p1 = {4{{4{(-2'sd1)}}}};
  localparam [5:0] p2 = (5'd2 * ((3'd7)^(2'd2)));
  localparam signed [3:0] p3 = {(~(((2'd0)<<(2'd0))?(2'd2):((4'd2)?(3'd4):(2'd0))))};
  localparam signed [4:0] p4 = (~^(4'd6));
  localparam signed [5:0] p5 = ((((-3'sd1)?(2'd2):(-3'sd1))/(2'd0))|(((5'd31)>(-5'sd11))<=((3'd1)>>(4'sd3))));
  localparam [3:0] p6 = ((4'd12)>>{((-4'sd2)?(-2'sd1):(3'd4))});
  localparam [4:0] p7 = ((|(~|(4'd1)))>=(2'sd0));
  localparam [5:0] p8 = (+((!(((2'd2)&&(5'd5))<<((5'd1)===(2'sd0))))&(~(^(((-3'sd0)<<<(3'd2))%(-3'sd3))))));
  localparam signed [3:0] p9 = (((^(+(-5'sd2)))>>{1{(3'd0)}})&&(+(^(((2'd2)>>(3'd2))>(+(5'd20))))));
  localparam signed [4:0] p10 = {{(4'd14)},(-(-5'sd13))};
  localparam signed [5:0] p11 = ((!((3'd1)||(3'd3)))%(-3'sd0));
  localparam [3:0] p12 = ({(2'd3),(5'd11),(-3'sd2)}-{(2'd2)});
  localparam [4:0] p13 = (|(4'sd1));
  localparam [5:0] p14 = ((((3'sd1)<<(4'd6))-{(4'sd2),(3'sd1),(3'd6)})+{2{(+(3'sd2))}});
  localparam signed [3:0] p15 = ((4'd14)!=(2'sd1));
  localparam signed [4:0] p16 = ((4'd6)?((5'd10)?(4'd3):(-4'sd2)):(3'sd1));
  localparam signed [5:0] p17 = (((4'd14)^((-4'sd0)%(4'sd1)))&&(-(~&((-4'sd3)?(5'd21):(3'd7)))));

  assign y0 = (2'd1);
  assign y1 = (((p3&&p14)&(~^p7))+({p13,p17,p4}&(a1?p10:p0)));
  assign y2 = ($signed((2'sd0))^~(5'd3));
  assign y3 = (6'd2 * (~(|p2)));
  assign y4 = (({2{(p8|p16)}}^{4{p3}})||(-({{a2,a5},(~a4)}!=={1{(a4<b4)}})));
  assign y5 = (({a2}|{b3,a4})!=={{2{b4}},(a3>>b2),(3'd3)});
  assign y6 = {(~|(^(&(3'sd2)))),(&{3{(p2>>>p8)}})};
  assign y7 = (({4{p6}})?$signed($unsigned({4{p10}})):$unsigned({3{p13}}));
  assign y8 = (-(~&$unsigned((b0>>a3))));
  assign y9 = (((b3!=b3)?(a0<p5):(a4&a4))>>((b1?a1:a0)?(b1&a4):(~&{a1,b1,p0})));
  assign y10 = (3'd5);
  assign y11 = {3{(p3<=p4)}};
  assign y12 = (((((b3>>>a3)<<<(p0|a3))-{2{{p12,b2,p11}}})|({{3{b0}},(a2<<<p14)}>>((a4|a2)<<<(a0&p0)))));
  assign y13 = (((a5&a4)<=(a5>>a4))<<(&(4'd2 * (~|{b0,a0,a1}))));
  assign y14 = ({(p10|p9),{b1,b5,a4}});
  assign y15 = ((+$unsigned(p1))?(p6&&p5):(|(-b5)));
  assign y16 = ($unsigned((($signed($signed((b2>a1)))^{{b1},(5'd2 * b2)})===$signed(({({($signed(a4))})})))));
  assign y17 = ((p10?p0:p3)?(p9?p9:p3):($signed(a5)<(p6?b4:b3)));
endmodule
