module expression_00912(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|((!(|{(((4'd1)==(3'd6))!==(~(-4'sd6)))}))>>>{(|(5'sd10)),(!(3'sd0)),((3'sd0)<<(4'd11))}));
  localparam [4:0] p1 = (-((|{2{{4{(5'd25)}}}})^~{4{(^(2'd0))}}));
  localparam [5:0] p2 = ({(3'd5)}<((-4'sd2)-(-5'sd9)));
  localparam signed [3:0] p3 = {{((-2'sd0)+(4'd11)),((2'd2)||(2'sd1))}};
  localparam signed [4:0] p4 = ((3'sd3)?(5'sd10):(2'd1));
  localparam signed [5:0] p5 = ((2'sd1)?(2'sd1):(4'd4));
  localparam [3:0] p6 = ((!(3'd0))-((3'd5)==((3'd4)?(2'd0):(4'd5))));
  localparam [4:0] p7 = (4'd2 * {1{((4'd6)>=(4'd4))}});
  localparam [5:0] p8 = {{(3'd3),(3'sd3),(2'sd0)},((-5'sd11)|(2'd1))};
  localparam signed [3:0] p9 = (~|(4'sd4));
  localparam signed [4:0] p10 = ({1{(-4'sd4)}}-(((3'd5)<(4'd2))>={1{(-3'sd0)}}));
  localparam signed [5:0] p11 = {4{{((-3'sd0)|(3'd4))}}};
  localparam [3:0] p12 = (3'd0);
  localparam [4:0] p13 = (-((-5'sd0)?(4'd6):(!(&(2'd3)))));
  localparam [5:0] p14 = (^{3{(~&(3'd7))}});
  localparam signed [3:0] p15 = ((5'd2)||((2'sd0)!==(-4'sd3)));
  localparam signed [4:0] p16 = (!((((5'sd11)?(5'sd7):(-2'sd1))/(4'sd1))>>(((5'd4)?(2'sd1):(4'sd3))%(3'd4))));
  localparam signed [5:0] p17 = ((((5'd20)-(4'd9))<<<{3{(-3'sd1)}})&({4{(-4'sd1)}}&((-4'sd5)===(5'd3))));

  assign y0 = $unsigned((2'd0));
  assign y1 = ((5'd18)==(~(3'sd2)));
  assign y2 = (^p3);
  assign y3 = ((|((a4?a5:a0)?(b3):{p9,b0,a0}))?$unsigned((4'd13)):((b2?b1:p2)?{4{p3}}:{1{b4}}));
  assign y4 = ({((p8||p14)^~(|p15)),(b1?a1:p6)}||(((p9^~p9)|(b5===b3))<=(~|(&(p1>=b1)))));
  assign y5 = (~(3'd5));
  assign y6 = (~(|(5'sd3)));
  assign y7 = {(({b0}-(b3>>p3))>($unsigned($unsigned({3{p0}})))),$unsigned({4{{1{p12}}}})};
  assign y8 = (-(-(4'd3)));
  assign y9 = {((p4?p3:a5)!=(p17?p1:p5)),(p7?p14:p9),(2'sd0)};
  assign y10 = ({3{(~|b0)}}?{1{(+((~^a2)<<<(a0)))}}:((a5?a3:a0)&&(-$unsigned(a1))));
  assign y11 = ($unsigned($signed((~&((3'd5)>(p7-p7)))))>>((b2+a5)%b0));
  assign y12 = {((4'd2 * p0)||{p9,p3}),({4{p13}}>>>{p10,a0,p13}),((p5&&p15)+(p17<<p10))};
  assign y13 = ({(a4?p0:p16),(p0!=p1),(~^p16)}&({a2,p13,a1}?{p11}:(b4|p16)));
  assign y14 = {{{1{{{3{a0}},{p12},(p13?p16:p11)}}}},{1{{2{(p7?b5:p2)}}}}};
  assign y15 = (|{{(&((p14&&b5)||(~^p4))),{{b1,p1},{p15,p9}},({a3,p11,a1}<{(~&b1)})}});
  assign y16 = (+(+(^(&((|(^(-(|(~|(!a5))))))>>>(~(~((^b4)!==(|b3)))))))));
  assign y17 = {(a4?a3:a4),(~&p16),(-a2)};
endmodule
