module expression_00763(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd11)?(-5'sd4):(3'sd1));
  localparam [4:0] p1 = {3{{2{{2{(5'sd8)}}}}}};
  localparam [5:0] p2 = {4{((-2'sd1)>=(-2'sd0))}};
  localparam signed [3:0] p3 = ((~|(-3'sd3))<((4'd14)|(5'd4)));
  localparam signed [4:0] p4 = (5'd1);
  localparam signed [5:0] p5 = {{(-{(2'd1),(4'sd5),(3'd2)})},(+{(3'sd1),(-5'sd2)}),{1{{(-5'sd6),(2'd2)}}}};
  localparam [3:0] p6 = {(-(^{(-2'sd0),(4'd10),(2'sd0)}))};
  localparam [4:0] p7 = (5'd2 * ((4'd13)-(3'd4)));
  localparam [5:0] p8 = {(!((-4'sd6)&(-5'sd7)))};
  localparam signed [3:0] p9 = (({(-3'sd3)}>={(-5'sd13)})&({(2'd1),(5'sd13),(5'd15)}===((-2'sd1)&(-3'sd1))));
  localparam signed [4:0] p10 = ((5'd30)?(2'd0):(2'sd0));
  localparam signed [5:0] p11 = (-3'sd2);
  localparam [3:0] p12 = (!{3{(((3'd6)==(4'd0))-(-(4'd8)))}});
  localparam [4:0] p13 = (((-5'sd14)|(2'd1))%(5'd1));
  localparam [5:0] p14 = (((4'd5)&&(2'sd1))<<(-4'sd5));
  localparam signed [3:0] p15 = ({3{{4{(-2'sd1)}}}}||(((2'sd0)&(-5'sd12))>>((5'd25)<<(-4'sd5))));
  localparam signed [4:0] p16 = (((~^(5'd11))?(^(4'd2)):{(3'sd0),(5'd3)})+{3{((4'sd1)?(2'd1):(3'd2))}});
  localparam signed [5:0] p17 = ({{(4'd6),(4'sd6),(3'sd0)},(~^{(-3'sd0),(4'd5)})}<<<{{((3'd5)|(5'd19)),{(3'd2),(3'sd1)},((-2'sd1)&(5'd3))}});

  assign y0 = $unsigned(a5);
  assign y1 = (-{1{b2}});
  assign y2 = {a2,a5,b4};
  assign y3 = ({(b4<=a0),{1{p3}}}>>({b5}^~(b1===a3)));
  assign y4 = $signed(a4);
  assign y5 = ((4'd13)^{(-2'sd1)});
  assign y6 = (((5'd2 * p6)-(p2-b0))!={{((b3-b3)!==(a1==b0))}});
  assign y7 = {(p7>=p13),(p4>p5),(p11<=b5)};
  assign y8 = (^(~&(~{(p14?p0:p5),{({a4})},(~{(~^p12)})})));
  assign y9 = {b4};
  assign y10 = ({4{a4}}?(b0?a4:b3):{4{a3}});
  assign y11 = (((b1?a0:a1)>(b4?a2:a0))>>({1{b5}}?$unsigned(a2):(a5^~b2)));
  assign y12 = {(b0?b0:b1),{{3{b1}}}};
  assign y13 = (|$unsigned((!(~|$signed((+$unsigned((!(^$unsigned($signed((^(~|(+(~|(&a3))))))))))))))));
  assign y14 = (+p12);
  assign y15 = (&(~&((a0>=b4)?(p1?a0:a5):(~^(b0===a1)))));
  assign y16 = ((p17?p12:b4)<<<(~|(+(-a1))));
  assign y17 = ({{p1,p16},(p7&&p5)}^~{{p15},(p16^~p15),(p8^~p8)});
endmodule
