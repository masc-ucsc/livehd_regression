module expression_00445(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd1);
  localparam [4:0] p1 = {4{{1{(5'd14)}}}};
  localparam [5:0] p2 = (((6'd2 * (3'd7))>>((3'd0)<(3'sd2)))<<<(((2'sd0)>>>(-2'sd0))-((2'sd0)>>(4'sd6))));
  localparam signed [3:0] p3 = (2'd2);
  localparam signed [4:0] p4 = (2'd0);
  localparam signed [5:0] p5 = (((4'd12)<=(5'd15))-((5'sd4)<<<(4'sd2)));
  localparam [3:0] p6 = (((5'd15)?(-5'sd3):(2'sd1))!=={1{(-2'sd0)}});
  localparam [4:0] p7 = (&{{(~(~^(!(|(~|(-4'sd4)))))),(+(|(!(~(~^(5'd16))))))}});
  localparam [5:0] p8 = (((5'sd3)<(2'd0))>>>(~^{(2'd2)}));
  localparam signed [3:0] p9 = ((-4'sd3)?(2'sd1):((2'sd0)?(3'd6):(-2'sd1)));
  localparam signed [4:0] p10 = {1{((!(5'd2 * ((4'd9)||(4'd15))))<={3{((2'd1)>>(-5'sd15))}})}};
  localparam signed [5:0] p11 = ((-5'sd12)^(2'd1));
  localparam [3:0] p12 = (|(4'd6));
  localparam [4:0] p13 = (~{{2{{((-5'sd4)==(-3'sd0)),((5'd20)-(-4'sd4))}}}});
  localparam [5:0] p14 = (2'd0);
  localparam signed [3:0] p15 = ((&({3{(3'sd2)}}&((-2'sd1)?(-2'sd0):(5'd24))))?(~&((~(-5'sd9))>>(-(5'd26)))):((~&(3'sd1))?{3{(4'd14)}}:(~&(4'sd2))));
  localparam signed [4:0] p16 = {{3{(5'd11)}},(^(3'sd2)),(((2'sd0)?(5'd8):(3'd4))==((-4'sd5)?(4'd2):(2'd3)))};
  localparam signed [5:0] p17 = ((((3'd2)/(-4'sd7))?((-3'sd3)<<<(3'sd1)):(-4'sd6))+(~(-(((3'd2)/(5'sd14))?(|(2'sd0)):((-4'sd2)?(-4'sd1):(2'sd1))))));

  assign y0 = ((~&((a3||b2)!=(a0?p6:a4)))||({2{b1}}?(b5!=a5):(a0?a1:a2)));
  assign y1 = ((((p11<p15)?(p17==a4):(a1+p1))>>((b1?a3:b3)?(p6?p10:p4):(b1?p12:a2)))<<<(((p14^a1)?(p17?a1:a0):(a4!==b3))<((p17|b1)^~(p7<<<b1))));
  assign y2 = (^((a1||a3)!=={a0,a5}));
  assign y3 = ({2{$unsigned((&(-($unsigned({1{{b2,b2,p4}}})))))}});
  assign y4 = (!a5);
  assign y5 = ((4'sd7)?(p8?a5:b1):$signed(p16));
  assign y6 = ({1{(b1?p13:a3)}}?((2'sd0)<=(p16>p15)):((4'sd0)==(p17>>a3)));
  assign y7 = (((5'd2)|(5'd29))||((5'd20)?(-2'sd1):(p5?p11:p5)));
  assign y8 = {(a2^~a3),{p11,b2},(b5<p16)};
  assign y9 = {1{(p11>=p16)}};
  assign y10 = (-(+{(~|(p12!=p13)),(p3==p3)}));
  assign y11 = (+($signed((!{2{(~^(~|a1))}}))^(((b3)>=(b3^~a4))!=={4{a3}})));
  assign y12 = (((~&a1)?(p14?p8:p11):(p0?p14:p16))?((p0?p3:p4)?(~&p4):(b2?b1:p2)):((^b1)?(+p1):(p14?p12:p6)));
  assign y13 = (-((+(^$unsigned({$unsigned({(b4),$unsigned(b0)}),((~(+$signed({b3,b5,b2}))))})))));
  assign y14 = (-3'sd3);
  assign y15 = {2{(&(|((b2|p1)<(a3?a1:p5))))}};
  assign y16 = ({4{(p1==p11)}}<=((p14>>>b5)||(p16==a0)));
  assign y17 = (p13||p2);
endmodule
