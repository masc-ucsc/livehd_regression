module expression_00923(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'sd1)?((-3'sd2)?(3'd3):(5'd27)):(2'd3))?(3'sd1):{((-5'sd8)?(5'sd15):(5'd14)),(6'd2 * (2'd3)),(4'd2)});
  localparam [4:0] p1 = {3{(((-3'sd2)?(-4'sd5):(5'd3))?{3{(5'd17)}}:{4{(5'd19)}})}};
  localparam [5:0] p2 = ((4'd5)===(5'd1));
  localparam signed [3:0] p3 = (-3'sd0);
  localparam signed [4:0] p4 = (~^{(-3'sd1),{1{(-2'sd1)}},(5'sd14)});
  localparam signed [5:0] p5 = {3{(-5'sd9)}};
  localparam [3:0] p6 = (-(4'd2));
  localparam [4:0] p7 = ((((4'sd1)>>(-4'sd2))>>{4{(-4'sd6)}})<=(-3'sd3));
  localparam [5:0] p8 = ((((5'sd2)!==(4'd4))?((3'd4)<=(3'd1)):{4{(4'd1)}})^~(2'd3));
  localparam signed [3:0] p9 = (((4'sd6)^~(5'd24))*(-(^(-2'sd0))));
  localparam signed [4:0] p10 = {4{(-5'sd5)}};
  localparam signed [5:0] p11 = {4{(2'd1)}};
  localparam [3:0] p12 = (-5'sd11);
  localparam [4:0] p13 = (~(5'sd0));
  localparam [5:0] p14 = (|(3'd0));
  localparam signed [3:0] p15 = (~&(2'd0));
  localparam signed [4:0] p16 = {4{(-2'sd1)}};
  localparam signed [5:0] p17 = (~{{((^((3'd0)===(3'd2)))!=={(2'sd0),(2'd1)}),{((2'sd1)+(4'd14)),{(3'd0),(5'd4),(2'd3)}}}});

  assign y0 = {{{4{{a5,p2,b5}}}}};
  assign y1 = {(~^(|(-{{(|(-(~|p4))),(&(4'd2 * p13))},((|(^(^p15)))>=(~(~(^p3))))})))};
  assign y2 = {3{{3{(2'd3)}}}};
  assign y3 = (4'd2 * {1{(p1==p2)}});
  assign y4 = (((b2!==b4)+(p14?b1:p6))>>(p15?b1:a2));
  assign y5 = (3'd6);
  assign y6 = {1{(|(~^(~|(({3{p16}}>>>(p11&p16))>>>((!p13)<<(p13>p0))))))}};
  assign y7 = {2{$signed((&(~&{p4,p6})))}};
  assign y8 = {(^(~&(2'sd1))),(^(~^(b0<<b2))),((a4>b5)!=={a1,a2,b0})};
  assign y9 = {1{(({2{(b2-b1)}}==$signed((p15^~a0)))|(({a5,a1,b4}>=(b0^~b0))>$unsigned((a2!==a5))))}};
  assign y10 = (~&((|(^{(a0<p8),{3{a1}},(b3<<<a5)}))>>({2{(p8>>a1)}}^{2{(b0-a5)}})));
  assign y11 = ((~^(+((b1)?(p17):(~&b1)))));
  assign y12 = (~&((!b2)));
  assign y13 = ((~^(&(|((b2<p1)>>(b3<a4)))))<<<(~((&(a2>>>a3))&(p13&&a4))));
  assign y14 = {(~^a4),(|p13),(~^p9)};
  assign y15 = ({({a2,a4,p12}?(p6!=p10):{2{a3}}),((p0&&p11)?(5'd2 * p8):(a1+b2)),{2{({p15,p11,a2})}}});
  assign y16 = {(a5>=p10),{(3'd0)},(a0>>>p6)};
  assign y17 = ((({p5,p12}>(b1+p8)))^({a2,b1,b3}>(+{b2,a5,b2})));
endmodule
