module expression_00233(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'sd0),(-2'sd0),(4'sd2)};
  localparam [4:0] p1 = ({3{(3'd2)}}?{4{(-2'sd1)}}:(2'sd0));
  localparam [5:0] p2 = {(|(~^(&(2'sd0)))),(3'd3)};
  localparam signed [3:0] p3 = (((!(4'sd3))?(+(4'd5)):{4{(5'd9)}})?{2{((5'd21)>(5'd20))}}:((~|(5'd18))||((-4'sd0)?(5'd23):(2'd1))));
  localparam signed [4:0] p4 = (6'd2 * {((5'd12)===(3'd3))});
  localparam signed [5:0] p5 = (-3'sd3);
  localparam [3:0] p6 = (((~{3{(-4'sd4)}})==(((5'sd13)==(3'd1))>={(-2'sd0),(-3'sd1),(4'd13)}))>({4{(-5'sd8)}}>{(|((2'd2)|(-4'sd0)))}));
  localparam [4:0] p7 = ((^(~|(((2'd1)|(-5'sd15))<<(4'd2 * (5'd26)))))!==((~((-3'sd2)^~(4'd0)))*((-3'sd0)<(2'd1))));
  localparam [5:0] p8 = (((4'd8)?(-5'sd0):(4'sd5))-((-4'sd4)||(4'sd2)));
  localparam signed [3:0] p9 = ((4'sd5)+((3'sd1)>>>(3'd5)));
  localparam signed [4:0] p10 = ({2{{2{(3'd1)}}}}<<(4'd0));
  localparam signed [5:0] p11 = (((3'd4)+(2'd3))%(3'd3));
  localparam [3:0] p12 = (~^(3'd4));
  localparam [4:0] p13 = ((4'd13)>=((((3'd0)&&(-3'sd3))^((2'sd0)>>>(5'd23)))&&(3'd6)));
  localparam [5:0] p14 = {{2{({{(4'd9),(5'sd12),(5'sd8)}}^{(|(5'd26))})}}};
  localparam signed [3:0] p15 = (2'd3);
  localparam signed [4:0] p16 = (3'd1);
  localparam signed [5:0] p17 = (~^(+(~(^(~^(|(+(!(+(~|(5'd25)))))))))));

  assign y0 = (|(~|((~&(+(a4?a2:b1)))?(a0?p12:b3):(a3?a2:a2))));
  assign y1 = (((b3/b2)^(b5?a0:b4))?((b1?b2:b2)==(b5*a5)):((a5?b4:a2)?(p11?b1:b3):(b4>>>a4)));
  assign y2 = {(3'sd1)};
  assign y3 = (-{4{(&p8)}});
  assign y4 = {(b2<=p0)};
  assign y5 = {3{((p6?p10:p15)>=(p14>>>p8))}};
  assign y6 = {({2{(p11>p7)}}),(4'd15)};
  assign y7 = (4'sd7);
  assign y8 = (((~$signed(b1))<<{p6,b5,b5})?(~((b3||a5)<=(-b2))):(~^{(&b1),(~&a2)}));
  assign y9 = ({((a5>a0)^~(p4>>>b1))}<=((a0?a0:b4)===(b2&&a2)));
  assign y10 = ((((~(p11+b0))&&$unsigned((p9<p16))))|((p12+a4)%p5));
  assign y11 = $unsigned((-(5'd11)));
  assign y12 = $unsigned({3{(~|p2)}});
  assign y13 = (((3'd5)<(2'sd0))||(-3'sd3));
  assign y14 = ((a4!==b2)?(a0>a5):(a4==b2));
  assign y15 = ($unsigned(((b1!==a3))));
  assign y16 = {((p7?p8:p8)^~(p15&p14))};
  assign y17 = (((((a5&a0)<={b1,a5})+(!((~|a3)))))===(((a4?b1:a2)-(~|b4))>={(b4?a5:a5)}));
endmodule
