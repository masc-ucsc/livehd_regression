module expression_00750(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-((~|((-2'sd0)!=(4'sd1)))!=((5'd26)||(-2'sd1))));
  localparam [4:0] p1 = (-(4'd14));
  localparam [5:0] p2 = (5'sd4);
  localparam signed [3:0] p3 = {4{(3'd4)}};
  localparam signed [4:0] p4 = ((5'd2 * {1{{(5'd27),(4'd13),(5'd1)}}})!==({(2'd0),(4'd11),(-5'sd15)}^~((3'd3)<<<(3'sd2))));
  localparam signed [5:0] p5 = (+(^({((-4'sd7)?(3'd3):(3'd7)),(~^(4'd15))}+{(2'd0),(2'd2)})));
  localparam [3:0] p6 = (5'sd0);
  localparam [4:0] p7 = ((3'd5)!=(-3'sd0));
  localparam [5:0] p8 = (-3'sd2);
  localparam signed [3:0] p9 = ({(2'sd0),(2'd2),(5'sd8)}^~{(-4'sd6),(3'sd0),(-3'sd2)});
  localparam signed [4:0] p10 = {(((4'sd4)>>(4'd5))>=((3'd4)|(5'd9))),(4'd2 * {(3'd1),(2'd0),(3'd5)})};
  localparam signed [5:0] p11 = ((-((4'sd3)>>>(2'd1)))!=(((3'd0)===(4'd7))<<((4'd8)>(2'sd0))));
  localparam [3:0] p12 = (((+(~(4'd6)))&&(-(~^(-2'sd1))))&(~^(~&({4{(2'sd1)}}===(~^(4'sd4))))));
  localparam [4:0] p13 = (({3{(2'd3)}}&&{(2'd3),(5'd29),(3'd3)})>={(~|(5'd3)),((2'd3)<=(5'd7)),((2'sd1)>=(3'd4))});
  localparam [5:0] p14 = ((+(5'd28))*(~(3'd5)));
  localparam signed [3:0] p15 = (((!(2'd0))?(+(-2'sd0)):((-2'sd1)?(2'd2):(4'd11)))?({(4'sd2)}?(-(3'd4)):{(-5'sd6),(5'd15)}):((&(-3'sd2))?((-4'sd7)?(-2'sd1):(4'd6)):((2'sd0)?(-4'sd0):(-3'sd0))));
  localparam signed [4:0] p16 = ((3'd7)>>((-2'sd0)!==(5'sd14)));
  localparam signed [5:0] p17 = (((!(-5'sd1))?((-3'sd1)?(2'd1):(-3'sd3)):((3'd2)?(-4'sd1):(4'd4)))>>>(((3'd0)/(4'sd2))?(|(2'd3)):(~|(-5'sd6))));

  assign y0 = (~&$unsigned(p11));
  assign y1 = $unsigned((($signed($signed(($unsigned($unsigned(($signed(($unsigned($unsigned($signed($signed((b1))))))))))))))));
  assign y2 = (~|(((5'd2 * (p6^~p8))>>((p8|p2)>=(b4-b3)))>>({1{(-(!a5))}}>>>((a4|p1)!=(a0!=b2)))));
  assign y3 = ((|((~^b5)>(b0<<a0)))|((b4>=b1)>(+(~a4))));
  assign y4 = {b4,p15,p4};
  assign y5 = (!p2);
  assign y6 = (4'd10);
  assign y7 = ((&{4{a4}})-((a1!=a5)&&(a0||a0)));
  assign y8 = (((5'd15)>=(a0?p1:a2))?((2'd0)<=(-5'sd7)):((a2?a3:b2)?(p14||p0):(a0!==a1)));
  assign y9 = {2{{3{(p7?p1:b4)}}}};
  assign y10 = {((~{p11,p12,p5})<<<(p4<<p15)),(~&((!(2'sd1))!=(p8|p9)))};
  assign y11 = (~^(~((~^((~^p7)>=(!p14)))^~(3'd1))));
  assign y12 = ((((a0&&b1)>>(!a1))>=((b4%a2)-(a0?b0:b4)))<<((3'sd2)?(b5||b2):(b0?a4:a3)));
  assign y13 = (&(~(~&{(!b3),(~&a4),{2{b0}}})));
  assign y14 = ({((p11?p11:a0)>>>((a1>>>b4)!==(b4?b2:a1)))}>=({p8,a1}?(p12+b0):(b5&&a1)));
  assign y15 = {3{(-2'sd1)}};
  assign y16 = (3'd3);
  assign y17 = (!{(a2===a2),{p2,p17}});
endmodule
