module expression_00690(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((&(~((-3'sd2)===(2'd0))))!=(4'd9));
  localparam [4:0] p1 = (((&((4'd5)?(5'd22):(3'd3)))&((3'd5)?(5'd24):(5'd28)))^~(((5'sd3)|(3'd7))&&(!(5'd2 * (3'd3)))));
  localparam [5:0] p2 = (((5'd5)>(5'd0))|((2'd0)|(-5'sd15)));
  localparam signed [3:0] p3 = (~^((5'd29)?(4'd15):(2'sd0)));
  localparam signed [4:0] p4 = ((^(&(&(4'sd7))))<(((2'd1)-(5'd21))<((4'd15)^~(2'd2))));
  localparam signed [5:0] p5 = (5'd22);
  localparam [3:0] p6 = (((4'd3)===(-4'sd3))-((5'd0)>>(-4'sd3)));
  localparam [4:0] p7 = (-((|((3'd1)>>(5'sd2)))!=(~^(-3'sd3))));
  localparam [5:0] p8 = ((|(~&(|(~^(+(-3'sd0))))))!=(-(+(3'sd2))));
  localparam signed [3:0] p9 = ((4'sd6)+{4{(4'd10)}});
  localparam signed [4:0] p10 = ((-((2'sd1)?(3'd7):(2'd0)))=={(+(&(5'd21)))});
  localparam signed [5:0] p11 = ((((-4'sd4)-(5'd23))-((5'd20)^~(-2'sd0)))!==(((2'd2)+(2'd3))^((3'sd1)==(2'd3))));
  localparam [3:0] p12 = (-4'sd5);
  localparam [4:0] p13 = (!(4'd0));
  localparam [5:0] p14 = (~^(+(|(~&(^(~|(~^(~^(!(~(-(~|(!(-(3'd1)))))))))))))));
  localparam signed [3:0] p15 = (5'sd11);
  localparam signed [4:0] p16 = {3{(2'sd0)}};
  localparam signed [5:0] p17 = ((((2'sd0)===(5'sd7))<<<{((3'd6)?(5'sd15):(4'sd6))})^{(~^(5'd16)),(~&(4'd7)),{(3'sd3)}});

  assign y0 = (-(~&((~&(|((~^a0)===(a1===a5))))>>>((b3+a3)!==(a4&a5)))));
  assign y1 = {(|((^p1)<(a2===a3))),((+(~p8))!=(p0<p3)),((p5^~p2)<(2'sd0))};
  assign y2 = {(~|(2'sd1))};
  assign y3 = ((p0?a0:b3)?(-4'sd2):(a1?b1:b2));
  assign y4 = (5'd6);
  assign y5 = {a0,p8,b5};
  assign y6 = ((2'd2));
  assign y7 = (3'd5);
  assign y8 = (|(^($signed((2'd3))||(|{1{(!(~^(&(~^(~&(3'sd3))))))}}))));
  assign y9 = ({b1,a2}==$signed({a1,a2}));
  assign y10 = (p9<<a4);
  assign y11 = $signed((a0*p3));
  assign y12 = {3{(b2>a3)}};
  assign y13 = (((p12>p17)^(p12^~p1))>{{p15},(b5===b5)});
  assign y14 = ($signed($unsigned($signed(({3{(p13?p10:p10)}})))));
  assign y15 = (3'sd0);
  assign y16 = {(!((-(~&((a3>b4)!==(b2<=a2))))!==(&{3{{3{a0}}}})))};
  assign y17 = {2{($signed($signed((b5&&p15)))^~(((b0)===(a0?a5:a2))))}};
endmodule
