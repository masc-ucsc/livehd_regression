module expression_00007(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-5'sd2);
  localparam [4:0] p1 = (|(~(+(~{2{(~((-2'sd1)+(5'd20)))}}))));
  localparam [5:0] p2 = ((4'd2)==(-2'sd0));
  localparam signed [3:0] p3 = (((4'd6)?(5'd6):(3'sd0))*(4'd2 * (2'd2)));
  localparam signed [4:0] p4 = ((((-4'sd3)-(3'sd3))?((-3'sd1)?(5'sd5):(2'd1)):((-3'sd0)?(3'd4):(2'sd1)))>>>(((3'd6)?(-5'sd9):(4'd1))^~(3'sd2)));
  localparam signed [5:0] p5 = (((4'd0)<<<(3'sd1))==((2'd3)&(4'sd4)));
  localparam [3:0] p6 = (({1{(4'sd1)}}?{4{(5'd28)}}:((-4'sd0)==(5'sd6)))===((|(2'd2))?(|(4'sd0)):((4'sd0)?(4'd12):(-4'sd6))));
  localparam [4:0] p7 = ((-2'sd0)!==(4'd5));
  localparam [5:0] p8 = {2{(6'd2 * ((3'd2)||(3'd1)))}};
  localparam signed [3:0] p9 = (3'd3);
  localparam signed [4:0] p10 = (({1{(2'sd0)}}>>>((2'sd0)>>>(4'd4)))>>>{2{((-5'sd15)>(3'd4))}});
  localparam signed [5:0] p11 = (+(-((4'd2 * (~&(|(2'd1))))!=(((5'd7)!==(2'd2))?(~(2'd1)):((5'd4)&&(2'd0))))));
  localparam [3:0] p12 = {1{(+(^(-(2'sd1))))}};
  localparam [4:0] p13 = (((3'sd1)!=((4'd13)>>>(3'd6)))<<<((5'd26)&(2'd1)));
  localparam [5:0] p14 = (!(4'd10));
  localparam signed [3:0] p15 = ((4'd2 * ((2'd2)!=(4'd11)))<<<(((5'sd0)!=(-2'sd0))!=(&((3'd1)<(4'sd6)))));
  localparam signed [4:0] p16 = (({(5'd15)}<((-3'sd0)&(-5'sd5)))^{(4'sd0),(3'sd0),(5'd14)});
  localparam signed [5:0] p17 = (!(4'd2 * ((3'd1)?(3'd3):(2'd1))));

  assign y0 = (((4'd5)^~(2'd3))?(-3'sd0):(b2?p7:p1));
  assign y1 = {(a1!=a1),{a2,b1}};
  assign y2 = ((((p6<<<p6)!=(a1!==b1))!=((p12>>b3)>(p12?p0:p3)))<<<{({p16}?(p7<p1):{3{p12}}),((p14||p10)>(p9&&p2))});
  assign y3 = (~^(2'd3));
  assign y4 = (p1+a1);
  assign y5 = (^({1{(4'd12)}}?((p12?p11:p1)&&(4'sd0)):(~^{3{(p8&p2)}})));
  assign y6 = {1{(({1{a0}}===(-4'sd5))!==(-5'sd9))}};
  assign y7 = (((b5===a0)&&$unsigned((a3*a3)))>>$unsigned(((a5^a1)>$signed(b1))));
  assign y8 = (^{{p17,p8},(p10<<p10),(-p6)});
  assign y9 = {$unsigned((5'd8))};
  assign y10 = (-2'sd1);
  assign y11 = (~&({(p15?a0:p10),(~|p11),(+p17)}?{(~|{(p14?p16:p9)})}:(~(|{(p6?b2:b3)}))));
  assign y12 = (~|$unsigned((~&{(3'sd3),(|(&(|{p4}))),$signed((+(|(p7&&p2))))})));
  assign y13 = {a0,p15,b3};
  assign y14 = (^(a3>p5));
  assign y15 = {3{b2}};
  assign y16 = {4{p7}};
  assign y17 = ({$signed((^{p9,p12}))});
endmodule
