module expression_00148(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~{3{((-2'sd0)?(4'd7):(-4'sd5))}})||{4{((2'sd0)===(3'd1))}});
  localparam [4:0] p1 = (+{{((~((-4'sd4)<(5'sd0)))&(~|((-3'sd1)!=(4'd2))))}});
  localparam [5:0] p2 = {4{{(4'd7),(3'd0)}}};
  localparam signed [3:0] p3 = ({4{((4'sd3)+(4'd3))}}+(4'd12));
  localparam signed [4:0] p4 = (|((-(+((2'd0)|(4'sd3))))<=(2'd1)));
  localparam signed [5:0] p5 = (|(3'sd0));
  localparam [3:0] p6 = (({(3'd6),(-5'sd1)}?((5'd6)||(2'sd1)):((-2'sd1)?(-5'sd1):(-4'sd7)))|(!{1{(~|(5'sd7))}}));
  localparam [4:0] p7 = (&(+(|(~|(&(~&(&(|(!(~&(-(+(~|(~|(+(3'sd1))))))))))))))));
  localparam [5:0] p8 = {3{(5'd27)}};
  localparam signed [3:0] p9 = (4'd1);
  localparam signed [4:0] p10 = ((~&(-5'sd15))<<<(~|(-(2'sd1))));
  localparam signed [5:0] p11 = (~|{(!((&(&(3'd5)))?(^(~&(3'd4))):((4'd6)==(5'd0))))});
  localparam [3:0] p12 = ((3'd5)?(3'd1):(4'd5));
  localparam [4:0] p13 = {(~^{(((4'd2)?(4'd11):(-3'sd0))?((-4'sd3)==(2'sd0)):((-5'sd13)>=(2'sd1)))}),(((-4'sd1)===(4'd9))|((3'd5)!=(2'sd1)))};
  localparam [5:0] p14 = {3{((4'd0)>(4'd11))}};
  localparam signed [3:0] p15 = ((5'd3)&((2'sd0)/(-5'sd2)));
  localparam signed [4:0] p16 = ((3'd5)&&(3'd3));
  localparam signed [5:0] p17 = ((((4'sd7)>>>(3'd7))^((2'd2)<=(-4'sd1)))>>(((4'sd7)==(2'sd0))||{3{(2'd2)}}));

  assign y0 = (((b5!=a0)!==(-2'sd0))!==((2'd2)^(b5>>b1)));
  assign y1 = (((a3?b3:a4)-(a0>>>p2))<({a4,p6,p17}||{2{p12}}));
  assign y2 = {3{(-3'sd3)}};
  assign y3 = $unsigned(({{3{(5'd5)}}}+({({a5}<<<(a1!==b1))})));
  assign y4 = {{(~|(~(-(((!(~^b1))^~(+{b5,b1,b3}))!={((~|a3)!={b5})}))))}};
  assign y5 = ((!p16)<<{a0,a1});
  assign y6 = ((3'sd3)*(5'd2 * p2));
  assign y7 = (3'd3);
  assign y8 = ((($unsigned((b0===a1))^{4{a3}})===(({1{a2}}<$signed(a4))>>>($signed(b3)>>>(a2^a5)))));
  assign y9 = (~((&(p0>a5))?(p0+p11):(p9?p2:p4)));
  assign y10 = {({b2,p16,b4}<=((b5<=a4)<<(b4|b3))),$unsigned(($signed(a4)?(p5==b1):$signed(b1)))};
  assign y11 = (((6'd2 * a1)==(a1%p1))+((b3/p6)!=(p10>p15)));
  assign y12 = ((({3{a2}}||((a5?b5:b1)))!=={(a1!=b2),(-b1),{b0,a0}}));
  assign y13 = (~$unsigned(((~&b3)^(-a5))));
  assign y14 = ((p15<p9)/p9);
  assign y15 = (~|(((p5?p5:p15))-((p3+p4))));
  assign y16 = ((2'sd1)<{{b0,p7,a5},({p5,a4,p2})});
  assign y17 = (-4'sd3);
endmodule
