module expression_00337(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^(&(-(^(+(~|(3'd6)))))));
  localparam [4:0] p1 = ((!{(3'd5),(-3'sd1)})?(~|((4'd3)?(4'd15):(4'sd2))):{(2'd2),(2'd0),(2'd3)});
  localparam [5:0] p2 = {2{{3{(2'd3)}}}};
  localparam signed [3:0] p3 = {3{(|((5'sd12)-(3'sd2)))}};
  localparam signed [4:0] p4 = (-4'sd3);
  localparam signed [5:0] p5 = (((4'd14)>=(-5'sd15))?((2'sd1)<(3'd1)):(~(-(3'd2))));
  localparam [3:0] p6 = (^{(2'sd1)});
  localparam [4:0] p7 = ({4{(-4'sd7)}}&&{2{(|(5'd14))}});
  localparam [5:0] p8 = (((&{4{(3'd0)}})>((5'sd14)+(-3'sd1)))^((^((2'd3)&(-5'sd6)))&(~(~(-4'sd4)))));
  localparam signed [3:0] p9 = (4'd10);
  localparam signed [4:0] p10 = ((3'd4)&&((!(+(5'd10)))<((-4'sd0)?(3'd2):(5'sd5))));
  localparam signed [5:0] p11 = {{(4'sd2),{(-2'sd0),(-5'sd0),(2'sd0)}},{3{(-4'sd7)}},{{4{(-5'sd8)}},(4'd13)}};
  localparam [3:0] p12 = (|(+(((+(5'd21))!=((5'd23)&(2'sd1)))!==(+((|(5'd18))||((4'd3)^(4'd3)))))));
  localparam [4:0] p13 = {3{{{1{{1{{1{(5'd14)}}}}}}}}};
  localparam [5:0] p14 = ((((5'sd1)*(2'd2))-((2'sd0)/(5'd9)))>>>(((5'sd8)>>>(4'sd5))||((2'd3)/(-5'sd9))));
  localparam signed [3:0] p15 = ((((-4'sd6)&&(4'd7))&((5'd26)<<(5'd6)))==((~((5'd12)%(4'd15)))%(4'd13)));
  localparam signed [4:0] p16 = ((-3'sd2)<=(2'd1));
  localparam signed [5:0] p17 = {1{(~(+(&({2{(5'd4)}}<<(~(!(4'd14)))))))}};

  assign y0 = ((a3?a2:a5)<$unsigned((a4>>a2)));
  assign y1 = {2{b4}};
  assign y2 = (p1<=p17);
  assign y3 = (!(^{{4{a3}},{(-5'sd9),(a0?a3:b3)},(~{3{a2}})}));
  assign y4 = (~^($signed((&(a5|a5)))<<<($unsigned(b0)>=(&b1))));
  assign y5 = (((b5|p3)?(p5):(p2?a0:b5))?((b3?a0:b4)?(p15?p10:p4):(a3?p5:b4)):((p15?p2:b0)?(p8?p15:p14):(p14||a2)));
  assign y6 = (3'd6);
  assign y7 = (~|(|((p16!=p6)>>>(p12&p0))));
  assign y8 = $signed($signed({$unsigned($unsigned({$signed(a0)})),((({a2}))),({a5,b4,a1})}));
  assign y9 = (~|(|({2{p10}}?(p11?p5:p0):(~(+p0)))));
  assign y10 = (({b2,b3,b5}==(~{a5,b5}))!==(|((b2-a3)+{a4,a2})));
  assign y11 = ((({a3,b3}>>>(a0^~a2))!=={2{(5'd2 * b2)}})^~{1{{2{(b2<<<a2)}}}});
  assign y12 = ($signed(a3)?(b3?b4:a4):(p10!=b5));
  assign y13 = (((b3&p1)>>>{1{(a3?p17:p7)}})&&{3{(b2<<p6)}});
  assign y14 = (!((p14?p6:a5)?(~(^(b1?b5:p2))):(p12?p9:a5)));
  assign y15 = (5'd11);
  assign y16 = (|{1{(4'd3)}});
  assign y17 = ((p8&p10)&(p11<p12));
endmodule
