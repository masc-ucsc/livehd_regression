module expression_00855(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd3);
  localparam [4:0] p1 = (^(!{(~|{(~^(2'd3)),((5'd9)^(4'd2)),((5'd14)==(2'd1))})}));
  localparam [5:0] p2 = ((~^{1{(4'd7)}})?{4{(3'sd0)}}:((-3'sd3)?(2'd1):(4'sd1)));
  localparam signed [3:0] p3 = (((+((4'd7)!=(3'd5)))!==(2'd0))<<((!((3'sd0)>=(-3'sd3)))>>>((2'd1)+(4'd3))));
  localparam signed [4:0] p4 = {((~^(5'd10))||((5'sd12)>>>(2'sd1)))};
  localparam signed [5:0] p5 = ((~&((^(2'sd1))<((5'd4)<=(2'd3))))===(!(-(~|(&((-2'sd1)<=(-4'sd7)))))));
  localparam [3:0] p6 = ((-5'sd12)|(-3'sd0));
  localparam [4:0] p7 = ((((3'd6)/(2'd2))!=(3'sd1))|((3'd7)!==(5'd21)));
  localparam [5:0] p8 = ((((-5'sd12)===(2'd1))<<((-2'sd1)|(4'sd3)))!=={((-2'sd0)&(4'd3)),{(3'd6)},(!(4'd15))});
  localparam signed [3:0] p9 = ((((-2'sd0)>=(-5'sd10))==((2'd2)&&(4'd6)))^(((-2'sd1)<<<(3'd4))===(-((5'd16)===(4'd6)))));
  localparam signed [4:0] p10 = (-(~(~(^(~&(&(~((-2'sd1)-(2'd1)))))))));
  localparam signed [5:0] p11 = {({((5'd12)&&(3'sd3)),((4'd10)<(4'sd4))}===(((5'd19)<<(5'd1))&&((-3'sd2)==(-5'sd9))))};
  localparam [3:0] p12 = ((5'd3)%(3'd4));
  localparam [4:0] p13 = {1{(|(+{4{(4'd13)}}))}};
  localparam [5:0] p14 = ((((3'sd3)!==(5'd31))!=((-3'sd1)<<(5'sd0)))>{1{(~^((-3'sd1)^~(5'sd4)))}});
  localparam signed [3:0] p15 = (4'sd7);
  localparam signed [4:0] p16 = ((-{(-4'sd2),(2'd3)})<{(^(3'd6)),((2'sd1)&&(-5'sd12)),((2'sd1)>=(-5'sd9))});
  localparam signed [5:0] p17 = ((~&((2'sd0)?(5'd25):(3'd4)))/(5'sd8));

  assign y0 = {3{{2{b1}}}};
  assign y1 = $signed(p12);
  assign y2 = ((~^(a5<b1))>>>(b3&b3));
  assign y3 = (~^({(&(3'd2)),$unsigned($signed(a0)),{1{{1{b0}}}}}<<<(4'd1)));
  assign y4 = (((&a3)<(p4<=p11))+(+{4{a0}}));
  assign y5 = (((5'sd14)?{4{p14}}:(p2?p8:p9))+{3{(-2'sd0)}});
  assign y6 = {{2{{1{b1}}}},((p15<=p14)>{4{b1}})};
  assign y7 = {2{(+{4{(5'd29)}})}};
  assign y8 = {((4'd14)?{{3{p13}},(~|p8)}:(4'sd2))};
  assign y9 = ((^((b5<<b3)===(b4!==b5)))<{((p4+p8)>>>(p16!=a0))});
  assign y10 = (p15&&p6);
  assign y11 = {1{(3'sd0)}};
  assign y12 = ((((~(~&b3))?(b2%b1):(b2&&p7))<<(((-a5)?(4'd2 * p8):(p2/p6)))));
  assign y13 = (((5'd17)-{2{(3'sd2)}})>=(((a3<=b2)&&(b1===b4))|(+(2'sd1))));
  assign y14 = (~^(~&(~&(+(((^p14)?(a0?p4:b1):(-p4))^(+(~^(-(~^(p13?p17:a4))))))))));
  assign y15 = ((4'd2 * (a0-p14))>{(a3-p11),{b2,b3,b4},{b4,p5,p10}});
  assign y16 = ({{{3{a5}}}}?({a5,a5,b5}||{1{(p11?a1:a5)}}):({3{a2}}-{2{a4}}));
  assign y17 = {3{(~({1{b2}}||(b0<=a2)))}};
endmodule
