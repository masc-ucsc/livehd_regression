module expression_00691(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'sd3)?(4'sd5):(-4'sd0));
  localparam [4:0] p1 = ((-2'sd1)/(-5'sd10));
  localparam [5:0] p2 = {4{(-5'sd11)}};
  localparam signed [3:0] p3 = (!(4'd2 * ((3'd0)/(2'd3))));
  localparam signed [4:0] p4 = ((((4'sd2)/(-5'sd12))/(5'd31))<<(~(|((^(-3'sd1))!=((5'd27)*(2'd1))))));
  localparam signed [5:0] p5 = (|(~(3'd1)));
  localparam [3:0] p6 = ((5'd2 * ((4'd14)+(2'd3)))+(+((2'sd1)^~((-5'sd5)+(5'sd2)))));
  localparam [4:0] p7 = (({((5'd19)<=(5'd26))}!=={(5'd21),(-3'sd3)})+{((-2'sd1)<=(5'd3)),(-(4'sd4)),{(2'd1),(4'sd7),(2'sd0)}});
  localparam [5:0] p8 = {{{{{(-2'sd0),(5'd29)}},(2'sd1)}}};
  localparam signed [3:0] p9 = (((2'sd0)?(-5'sd9):(-2'sd0))?((3'd4)?(2'd0):(2'sd0)):((3'sd2)?(3'd5):(3'sd0)));
  localparam signed [4:0] p10 = (3'd1);
  localparam signed [5:0] p11 = ({1{((4'd0)?(3'd1):(3'd3))}}?((5'd30)-(-5'sd7)):((4'd1)>=(5'sd8)));
  localparam [3:0] p12 = ((5'd11)<(-3'sd2));
  localparam [4:0] p13 = (!(3'sd0));
  localparam [5:0] p14 = ((5'sd7)>>(-3'sd0));
  localparam signed [3:0] p15 = {(5'd16),(5'sd0),(3'sd2)};
  localparam signed [4:0] p16 = (!(4'd3));
  localparam signed [5:0] p17 = (((-2'sd1)===(3'd0))!==(&(&(3'sd1))));

  assign y0 = (2'd1);
  assign y1 = $signed(((((|b0)===(^b5)))>>>(~|((p11^~p1)/p3))));
  assign y2 = (4'd1);
  assign y3 = ({{p9,p0},{p5,p1},((p1-a1))}<=(-4'sd1));
  assign y4 = (((p7?p7:p4)>=(p13!=p2))<<({(p5^p2)}||(p0?p7:p11)));
  assign y5 = (~^(^{(+(a5?p1:a3))}));
  assign y6 = (~&(((&p0)>>>(p10<<<a0))^~((p0>>p2)<<$unsigned(p7))));
  assign y7 = {{(-5'sd11)},(~(|{(^a0),{b3,p14},{1{a1}}}))};
  assign y8 = ((+a1)!=={a4,b2});
  assign y9 = ((p9<<p3)?(b1!==b0):{p15});
  assign y10 = {4{(b4>>b2)}};
  assign y11 = {(+(p5&&a4)),((p17==p10)&&{3{p13}})};
  assign y12 = {{((b5&b1)>>(5'sd4))},{{{p12,p17,p17},(4'd8)}}};
  assign y13 = {{(a1+p4)},((p5||p6)|{a4})};
  assign y14 = {(-5'sd9),{(b5?b4:b3)},(a3?a4:b1)};
  assign y15 = (~{(!(^p1)),{(^p13)},{(^p17)}});
  assign y16 = (2'd1);
  assign y17 = ((b0==p7)>={1{p3}});
endmodule
