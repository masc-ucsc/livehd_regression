module expression_00965(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+((^{{(2'sd0),(4'sd1)}})?{(-4'sd3),(5'd25),(2'd3)}:((-2'sd1)?(4'd0):(-3'sd1))));
  localparam [4:0] p1 = (+{(2'd3),(3'sd1),(2'd2)});
  localparam [5:0] p2 = (+(~(2'sd0)));
  localparam signed [3:0] p3 = (((2'd2)?(4'd5):(5'd11))<((2'd1)||(3'sd3)));
  localparam signed [4:0] p4 = (({(3'd7),(4'd6),(2'd1)}!=((5'd24)?(4'd13):(2'd1)))?{((4'sd2)^(3'd0)),((-2'sd0)?(2'd1):(3'd7))}:({(4'd6)}<(&(-5'sd3))));
  localparam signed [5:0] p5 = (2'd2);
  localparam [3:0] p6 = (+(-((-5'sd0)?(5'sd7):(5'sd5))));
  localparam [4:0] p7 = (6'd2 * (4'd5));
  localparam [5:0] p8 = (((-4'sd3)>(3'd0))===(5'd30));
  localparam signed [3:0] p9 = ({(4'd12),(|(2'd0)),{(2'sd1),(3'd5)}}?{(-3'sd0)}:(((2'd2)?(-5'sd10):(2'sd1))<<<((5'd13)?(5'sd3):(-3'sd1))));
  localparam signed [4:0] p10 = ({1{(&((-5'sd8)?(-4'sd1):(3'd4)))}}||((2'd2)<<<((4'd2)!=(4'd11))));
  localparam signed [5:0] p11 = {4{{3{(4'sd7)}}}};
  localparam [3:0] p12 = ((~&(5'd12))?((4'd5)?(4'd7):(4'sd7)):((-3'sd2)?(-5'sd5):(-5'sd9)));
  localparam [4:0] p13 = {2{{3{((4'd5)||(3'sd1))}}}};
  localparam [5:0] p14 = {((2'd0)>>>(5'sd4)),(~(-5'sd3)),(~|(-2'sd1))};
  localparam signed [3:0] p15 = (4'd10);
  localparam signed [4:0] p16 = (4'd12);
  localparam signed [5:0] p17 = ((2'd2)^~(-4'sd1));

  assign y0 = (~^{((5'd28)^{(4'd11),(p1&&p15)})});
  assign y1 = (~&{3{{3{(+a3)}}}});
  assign y2 = (~|(((~^(a1>p1))?(p3!=p9):(p15^~p11))&(&(-(~(~((p3<<p11)/p14)))))));
  assign y3 = $unsigned(({(~^(p13>>>p2))}+({p7,p8,p16}!=$unsigned(a5))));
  assign y4 = (3'sd0);
  assign y5 = ({4{(b5>a2)}}||$unsigned($unsigned({1{((a4<b2)-(b4!==a3))}})));
  assign y6 = (+p12);
  assign y7 = (^(-(5'd8)));
  assign y8 = (+($unsigned((!(((-$signed(p17))?(a4?p9:b0):(+(^a5))))))));
  assign y9 = {(3'sd2)};
  assign y10 = ((b0?b4:a2)^~{p16,a5});
  assign y11 = (|a3);
  assign y12 = {({(p2?p14:p5)}<=(p17>p8)),(3'sd0)};
  assign y13 = {3{a0}};
  assign y14 = (-5'sd0);
  assign y15 = (-4'sd0);
  assign y16 = ((2'd1));
  assign y17 = ((((a3>>p7)+(^a0))<<((&p5)>={p4,p11}))>({(b1===b3),(p1<<<b5)}<<(^(!(a5&b2)))));
endmodule
