module expression_00403(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-5'sd14)?{4{(5'sd6)}}:(5'd17));
  localparam [4:0] p1 = ({(3'sd3),(5'd11),(5'd21)}^{(4'sd0)});
  localparam [5:0] p2 = ((~&(+{2{(2'd2)}}))||{2{{3{(3'sd2)}}}});
  localparam signed [3:0] p3 = ((4'd3)>(-5'sd6));
  localparam signed [4:0] p4 = {4{(4'd14)}};
  localparam signed [5:0] p5 = ((~|(~&((4'd1)?(4'd13):(5'd25))))<=(((4'sd2)+(4'sd2))===((2'd2)?(5'sd0):(5'd19))));
  localparam [3:0] p6 = (+(-(({1{(3'd5)}}===(~^(3'd2)))!=(!(~&(!(~|(-3'sd3))))))));
  localparam [4:0] p7 = ((((-4'sd0)||(2'sd0))<=((2'sd0)/(2'd3)))&&(((2'd2)===(4'd2))%(2'sd1)));
  localparam [5:0] p8 = ((!{1{(((-4'sd3)^~(5'd0))<(|(-4'sd1)))}})<<<({2{(2'd2)}}?((3'd7)?(5'sd15):(2'sd1)):{(4'sd1)}));
  localparam signed [3:0] p9 = ((5'd2 * (~^((2'd1)<<(3'd3))))>=(~^(-{3{(-5'sd14)}})));
  localparam signed [4:0] p10 = ((((5'd28)!==(2'sd1))>=(5'd12))<<<((5'd2 * (4'd12))!=((5'sd3)>>>(5'd31))));
  localparam signed [5:0] p11 = {4{(~&(3'd1))}};
  localparam [3:0] p12 = (((2'd1)+(-5'sd13))?((3'sd1)?(-5'sd9):(5'd30)):{4{(3'd3)}});
  localparam [4:0] p13 = ((((2'sd0)|(4'sd6))?((2'sd0)+(2'd1)):((-4'sd3)<<<(2'd0)))^(((2'sd1)!==(-3'sd1))+(4'd4)));
  localparam [5:0] p14 = (((-2'sd1)==(2'd3))*((4'sd2)!==(3'd1)));
  localparam signed [3:0] p15 = ((3'd4)<(2'd0));
  localparam signed [4:0] p16 = (((-3'sd1)<<<(5'sd0))>((5'd15)<(5'sd2)));
  localparam signed [5:0] p17 = ((-5'sd3)|(4'sd2));

  assign y0 = (~^(~^((b2%b5)|(~^(~^p13)))));
  assign y1 = ((b3!=b2)!==(b2|a2));
  assign y2 = $signed(((+{$signed(((^b0)>>$signed(a1)))})));
  assign y3 = (a3^p15);
  assign y4 = (5'sd0);
  assign y5 = $unsigned($unsigned(($signed(a3)<<<$unsigned(b4))));
  assign y6 = (-((-(a2>a2))));
  assign y7 = (((-5'sd6)===(5'd24))|(-5'sd9));
  assign y8 = {1{{3{{2{(p6&&p9)}}}}}};
  assign y9 = {4{{b1,b2}}};
  assign y10 = {{{2{(^{3{b5}})}},{1{{(~|(p9+b0)),(4'd2)}}}}};
  assign y11 = ((p17|p1)||(^(p12==p11)));
  assign y12 = ((2'sd0)^~((~^(p17?p6:p7))>>((p14>>>p17)<=(2'd0))));
  assign y13 = (|(^((+(&$signed(($unsigned($unsigned(p2))&(p14*b1)))))||(-(~^($unsigned((b0))<=$signed($signed(a5))))))));
  assign y14 = {3{(~&a4)}};
  assign y15 = ({b2,a3,a1}&(-(~(|b3))));
  assign y16 = (~^((!a1)?(b5<<<b2):$signed(p11)));
  assign y17 = ((p9&&p3)?{a5}:(5'd2 * b2));
endmodule
