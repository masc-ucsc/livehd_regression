module expression_00820(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(|(3'sd2)));
  localparam [4:0] p1 = {((3'sd1)-(-3'sd2)),((4'd6)!==(3'sd3)),(-(-4'sd2))};
  localparam [5:0] p2 = (((-2'sd0)^(-2'sd1))>>((4'sd2)?(2'd0):(4'd3)));
  localparam signed [3:0] p3 = ((~&{4{(3'd3)}})==={((-3'sd0)==(3'd3))});
  localparam signed [4:0] p4 = ((-2'sd0)===(+(~&({(2'd0),(2'd3),(4'sd0)}>(4'd1)))));
  localparam signed [5:0] p5 = {((4'sd0)+(-4'sd2)),((-3'sd2)<<(-2'sd0)),{(5'd7),(-2'sd1)}};
  localparam [3:0] p6 = (({4{(4'd4)}}||((-4'sd2)>>>(3'd0)))&{1{(-(^{4{(2'd3)}}))}});
  localparam [4:0] p7 = (((-3'sd0)&&(5'd4))&((2'sd0)?(2'd2):(2'sd1)));
  localparam [5:0] p8 = (((2'd0)^(4'd4))>>>(&(3'd2)));
  localparam signed [3:0] p9 = (!(~&(!(~(~|(~|(^(~&(&(^(|(~|(~^(^(-4'sd4)))))))))))))));
  localparam signed [4:0] p10 = (-(((4'd7)<=(^(5'd24)))&(-2'sd0)));
  localparam signed [5:0] p11 = {1{{1{((5'd8)?(4'd4):(4'd10))}}}};
  localparam [3:0] p12 = (-{(4'sd5),(3'd0),(3'sd3)});
  localparam [4:0] p13 = {(5'sd5),(5'sd14)};
  localparam [5:0] p14 = (2'd0);
  localparam signed [3:0] p15 = (^(+{1{{4{{3{(-2'sd1)}}}}}}));
  localparam signed [4:0] p16 = ((((3'd6)===(3'sd3))&{(-2'sd1)})>>(((-5'sd9)===(5'd4))>=((2'sd1)<(4'sd5))));
  localparam signed [5:0] p17 = (|(((~|(4'd15))>>((5'd14)!==(5'sd11)))?(-((-5'sd4)?(-3'sd0):(3'sd1))):(&((&(-5'sd8))===(&(4'd15))))));

  assign y0 = ((|(b2>=b0))!==(~|(&(&b1))));
  assign y1 = {1{(|(+p4))}};
  assign y2 = ((((!a3)===(a2-b1))>>(~(b2||a1)))&&(~&((+(p5^~p10))>>>(b2?p14:p15))));
  assign y3 = ((!((a4&&b4)===(a1<=b3)))^((p6>>p15)-(~p4)));
  assign y4 = (((a3!==b4)*(~&p10))<<<(~|(3'd3)));
  assign y5 = ((2'd0)==(3'sd3));
  assign y6 = (&(3'd7));
  assign y7 = (!(^{4{(-(~p17))}}));
  assign y8 = ((2'd2));
  assign y9 = (b5?p5:b3);
  assign y10 = $unsigned($unsigned(((($signed(p8))))));
  assign y11 = {(^{2{$signed(p14)}}),{(-(^{1{p5}}))}};
  assign y12 = (({p6,p9,a2}>={3{p5}})+((b5!==a3)==(b2!==a3)));
  assign y13 = {b3,b1,b3};
  assign y14 = (+(^$signed((6'd2 * (~|(-p1))))));
  assign y15 = (((4'd2 * (4'd4))^{2{(p11&p1)}})>=(((4'd3)!=(b0|b4))<=(-(p7<<p0))));
  assign y16 = ({(a4?a4:p3),(~p3)}?{4{b0}}:(3'd1));
  assign y17 = (!((p2?p13:p9)>>>(b5!==a2)));
endmodule
