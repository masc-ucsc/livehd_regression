module expression_00776(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-(4'd6))>=((2'd0)^(2'd1)));
  localparam [4:0] p1 = ((((3'sd1)!=(2'sd0))||{(-3'sd2)})+((5'd24)?(3'sd0):(-2'sd0)));
  localparam [5:0] p2 = {(((2'd2)?(3'sd2):(5'sd6))?{(5'd14),(5'd21)}:(~|(-3'sd2))),({(5'd17)}?(~(2'd3)):(&(-3'sd0)))};
  localparam signed [3:0] p3 = ((+(((2'sd0)>(-5'sd2))<<{(5'd27),(-2'sd0),(-5'sd10)}))!==(~&{(-(!(~^(-2'sd0))))}));
  localparam signed [4:0] p4 = {{(^{((5'd1)^~((3'sd1)===(5'd8))),(~^((3'd6)?(2'd1):(-4'sd5)))})}};
  localparam signed [5:0] p5 = {1{(((3'd4)^(2'd0))<((2'd3)<<<(4'd14)))}};
  localparam [3:0] p6 = {4{((5'd11)?(4'd4):(4'd0))}};
  localparam [4:0] p7 = {4{(-4'sd4)}};
  localparam [5:0] p8 = ((-2'sd1)?(4'sd7):(-2'sd0));
  localparam signed [3:0] p9 = (((5'd21)&(-5'sd11))?((3'd2)?(-3'sd2):(-5'sd7)):(~^(5'sd0)));
  localparam signed [4:0] p10 = {4{((3'd1)+(-4'sd2))}};
  localparam signed [5:0] p11 = (-(~|(+(~|(~(-(|(|(&(2'd3))))))))));
  localparam [3:0] p12 = (2'd1);
  localparam [4:0] p13 = (5'sd1);
  localparam [5:0] p14 = ((3'd0)?(-3'sd0):(-4'sd2));
  localparam signed [3:0] p15 = ((5'd15)<<(5'd23));
  localparam signed [4:0] p16 = ((~(-(~^((3'sd1)<=(2'sd1)))))&&(|(~|(~&((3'd5)||(3'sd1))))));
  localparam signed [5:0] p17 = (5'd2 * ((3'd1)-(2'd3)));

  assign y0 = $unsigned((((!p12)<(p9<=a5))>>$signed((^(p10|b2)))));
  assign y1 = (a4>p10);
  assign y2 = $signed({p4,p3});
  assign y3 = (!{{((6'd2 * {3{p12}})<(&({4{a3}}||(p4||b2))))}});
  assign y4 = (((((p5*p7)))<<<((p10^~p0)))==($unsigned((b3%b0))-$signed((p7<<<p16))));
  assign y5 = (b5<a1);
  assign y6 = ((b3&&b5)>=(p7^b5));
  assign y7 = (~^(((p16<<b0)<<<(a1|b0))&((a5==a1)!==($signed(a0)))));
  assign y8 = {1{((~^{1{(p16?p13:p5)}})&&((b4&p1)?(p15-a3):(p9>>p2)))}};
  assign y9 = {($unsigned(((p0==p7)<<{b1}))||$unsigned(((p4>>>p8)<(p13?p16:p12))))};
  assign y10 = (~^(-4'sd3));
  assign y11 = {4{{1{(5'd8)}}}};
  assign y12 = {(~^$unsigned((&{a4,p12}))),{{1{p2}},(-a4)},$signed({(-(p14))})};
  assign y13 = {p11,p13,p13};
  assign y14 = {{(~&{3{p12}}),{1{{p11,p4}}},(2'd1)}};
  assign y15 = ((b2&&a1)!=(b0&a0));
  assign y16 = (($signed($signed(b0))>(a2?p2:b3))?((-5'sd10)?$unsigned(a2):(3'sd1)):(3'sd3));
  assign y17 = (~&(~^{{{a1}},{b0,b3,b5}}));
endmodule
