module expression_00019(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd2);
  localparam [4:0] p1 = {{3{((2'd2)>>>(-5'sd3))}},{{(3'd1),(4'd10)},{4{(4'sd3)}},{(2'sd0),(3'd2)}}};
  localparam [5:0] p2 = (((-5'sd11)===(-5'sd0))||(~&((4'd4)?(3'd3):(-2'sd0))));
  localparam signed [3:0] p3 = {3{(5'd25)}};
  localparam signed [4:0] p4 = ((((5'd14)|(3'd1))!={(5'd15),(3'd3),(4'sd3)})||{((5'sd11)!=(4'sd6))});
  localparam signed [5:0] p5 = (5'd2);
  localparam [3:0] p6 = (-{1{(+((~^(2'sd1))<<{1{(3'd1)}}))}});
  localparam [4:0] p7 = ((^(6'd2 * (3'd1)))^~((&(-4'sd6))<(~|(-2'sd1))));
  localparam [5:0] p8 = ((2'd0)>>(5'd0));
  localparam signed [3:0] p9 = (((~&(5'd6))&&(4'sd5))?{3{((3'd4)>=(5'd17))}}:((5'd2 * (3'd0))?(6'd2 * (5'd18)):((-4'sd0)<<(3'd5))));
  localparam signed [4:0] p10 = {1{(3'sd2)}};
  localparam signed [5:0] p11 = ((5'sd13)<(2'd1));
  localparam [3:0] p12 = {(2'd2),(2'd0),(5'sd6)};
  localparam [4:0] p13 = ((2'd1)?(5'sd2):(4'sd6));
  localparam [5:0] p14 = {1{(+(~&(-3'sd3)))}};
  localparam signed [3:0] p15 = ((((+(2'd3))+(~&(-4'sd6)))-(|((3'd1)?(2'd3):(2'sd1))))-(!{3{((5'd28)!=(3'd1))}}));
  localparam signed [4:0] p16 = {4{(~^(3'd0))}};
  localparam signed [5:0] p17 = (2'sd0);

  assign y0 = (2'd2);
  assign y1 = (-((-{1{((p2||p17)^~(p7-p12))}})>>$unsigned($unsigned({3{{p5}}}))));
  assign y2 = (~^(((p15==p6)-(b1<<p4))<<((p8<=p14)|(a0<<<p2))));
  assign y3 = ({({a1,a4,a1}),(|(|b0)),((b4))}===$unsigned({3{(a2>>>b3)}}));
  assign y4 = {({(b2^~a0),(-(5'd2 * b1)),{1{(5'd16)}}}=={((4'd12)-{4{a3}})})};
  assign y5 = (~^(($signed((~(b2&b0))))!==({1{a3}}==(|b4))));
  assign y6 = $signed((~&($signed((~|(&$unsigned((+(p8&p17))))))||(((b1&b0))===((a2<b4)<=(a3==a3))))));
  assign y7 = $signed((!(+(-4'sd3))));
  assign y8 = {3{{{2{(|p6)}}}}};
  assign y9 = ((!(p3))|(4'd2 * p14));
  assign y10 = {b4,b1,p12};
  assign y11 = $signed($unsigned(p11));
  assign y12 = {a0,a1,p0};
  assign y13 = ((~&((p7?p3:p1)?(-a1):$unsigned(p14)))?(|(((~p2)?(|p3):(a3?p6:p1)))):((p2?p13:a5)?(~|p7):(p5?p5:b2)));
  assign y14 = {1{(&(^$signed(($signed((~|(^a3)))))))}};
  assign y15 = ((~^({4{a3}}>=((a1>p14)<(b0>b3))))||(((b4+b4)^(b3+a3))!==(!((a5^~a4)>=(a3&b5)))));
  assign y16 = (^(~|(-(~^(3'sd2)))));
  assign y17 = (((&(p4||a0))?(p8/p1):(b3|a0))+(+(&(~(~&(~&(b2?a5:p4)))))));
endmodule
