module expression_00036(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(((!(+(3'sd2)))&((-3'sd2)+(-4'sd4)))&&((~^(|(-2'sd1)))-((3'sd3)>>>(5'd6)))));
  localparam [4:0] p1 = (((4'd9)>(4'd0))<<(2'd2));
  localparam [5:0] p2 = (((~&(2'sd0))?((3'sd2)?(3'sd2):(-2'sd0)):((-5'sd3)!=(3'd5)))+{2{(|((5'sd5)?(4'sd4):(3'd5)))}});
  localparam signed [3:0] p3 = {4{((-3'sd2)?(5'sd11):(4'sd4))}};
  localparam signed [4:0] p4 = {4{(~|(-4'sd1))}};
  localparam signed [5:0] p5 = ((((-5'sd2)?(2'd3):(-4'sd1))?(2'd2):((5'd30)?(2'sd1):(-4'sd6)))|(4'd5));
  localparam [3:0] p6 = ((&({(-3'sd1),(3'sd3),(4'sd5)}<<<{4{(3'sd0)}}))!==((+(3'd3))?(&(-4'sd0)):((2'd1)===(4'd9))));
  localparam [4:0] p7 = (-3'sd2);
  localparam [5:0] p8 = (((2'd0)<=(3'd4))/(5'd21));
  localparam signed [3:0] p9 = (~|((((2'd1)>(2'sd1))?((2'd2)>>>(4'sd7)):{1{(-4'sd6)}})!=={1{(~|(~{2{((2'd3)?(2'd0):(4'sd4))}}))}}));
  localparam signed [4:0] p10 = (((~&(3'sd3))?{(4'sd3)}:{2{(2'sd1)}})^~(((-5'sd1)?(2'd1):(5'd29))<{1{(^(3'sd1))}}));
  localparam signed [5:0] p11 = (5'd2 * ((4'd11)>>>(5'd21)));
  localparam [3:0] p12 = {3{(5'sd8)}};
  localparam [4:0] p13 = {2{{((6'd2 * (2'd0))^~{4{(3'sd1)}})}}};
  localparam [5:0] p14 = {2{((~^((2'sd1)||(4'd9)))^{(-5'sd0),(4'd6)})}};
  localparam signed [3:0] p15 = ({{{(5'sd3)},((4'd0)+(3'sd1)),((3'sd0)<(-2'sd1))}}!=={((-3'sd0)^(3'd2)),((-3'sd0)||(-2'sd0)),((-3'sd1)-(5'sd0))});
  localparam signed [4:0] p16 = (((-4'sd2)?(5'd11):(5'd14))||(((3'sd2)<<<(2'd0))>>>(~(2'd3))));
  localparam signed [5:0] p17 = ((|{3{(-5'sd3)}})+(+((3'd3)|(2'sd0))));

  assign y0 = {(+($signed(b3)?(-p16):(-a0))),((p8?a2:b2)?(^b0):{p8,b1})};
  assign y1 = {1{($signed($signed({2{$unsigned((b3!==a3))}}))!==$signed($unsigned({3{{4{a1}}}})))}};
  assign y2 = (~p11);
  assign y3 = {(3'sd3),({p10,p7,p8}>={p17}),{4{a3}}};
  assign y4 = $signed(($signed(({3{b1}}>{4{b0}}))-{((b0&b2)),$unsigned((b1+a0)),$signed((a1|b3))}));
  assign y5 = {3{(a0===a0)}};
  assign y6 = ((-(-5'sd14))?$signed({1{{3{p16}}}}):($signed(a0)==={b5,a3,a2}));
  assign y7 = ((~|((b2<=p14)==(a3!=b0)))+(-((~&(a4*a0))===(4'sd5))));
  assign y8 = (|(-$signed({2{(3'd3)}})));
  assign y9 = (~^{4{(~{4{a1}})}});
  assign y10 = ((2'd2)?((b3<p2)^{p13,p4,p0}):({2{p12}}|(p17-b5)));
  assign y11 = {2{{3{(-3'sd0)}}}};
  assign y12 = {4{(b1||a5)}};
  assign y13 = ((((a0?p7:a2)^{4{a0}})>=((b1?a1:b1)<<(b3>a3)))>>((4'd2 * b2)?{2{b4}}:(b1>b4)));
  assign y14 = ((-2'sd1)?$unsigned((4'd8)):($signed(p13)?(-2'sd0):(b3===b1)));
  assign y15 = (~b5);
  assign y16 = ((-5'sd13)+(p4?p5:p0));
  assign y17 = (({p13,p5,p12}<<<(!p16))<<<(3'd1));
endmodule
