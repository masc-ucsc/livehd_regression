module expression_00542(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-((~|{1{(-2'sd0)}})>>>(^((-5'sd2)?(5'sd6):(-5'sd9)))));
  localparam [4:0] p1 = (&(4'd6));
  localparam [5:0] p2 = {3{(((-3'sd3)>=(5'sd5))+((-5'sd15)!=(5'd27)))}};
  localparam signed [3:0] p3 = ((-(6'd2 * (3'd5)))>((5'd13)!==(3'sd3)));
  localparam signed [4:0] p4 = {(5'd2 * ((3'd1)?(4'd1):(2'd0))),(+{4{((2'd3)?(-4'sd2):(2'sd1))}})};
  localparam signed [5:0] p5 = (((^((4'sd1)>>(5'd0)))<=((-(5'sd7))>((2'd2)>=(-4'sd1))))+(((!(4'sd3))>=(6'd2 * (4'd4)))|(2'd0)));
  localparam [3:0] p6 = ((-3'sd2)<((2'sd1)?{2{(-3'sd1)}}:((2'd2)?(3'd1):(2'sd0))));
  localparam [4:0] p7 = {3{(~&(-4'sd3))}};
  localparam [5:0] p8 = (^(&(((3'd5)<=(2'd1))^~{1{(3'd1)}})));
  localparam signed [3:0] p9 = (((3'sd0)===(3'sd2))!==((5'd20)<<<(3'd3)));
  localparam signed [4:0] p10 = (3'sd1);
  localparam signed [5:0] p11 = (((-4'sd5)^~(5'd15))>>>(((4'd4)||(3'sd1))>((-5'sd8)&(-2'sd0))));
  localparam [3:0] p12 = (((2'sd1)^(-4'sd6))?(2'sd0):((4'sd4)&(5'd2)));
  localparam [4:0] p13 = ((((2'd2)+(4'sd2))&&(+(~|(5'd4))))<<<(&((2'd0)^~(-(5'sd1)))));
  localparam [5:0] p14 = (((4'sd4)+(5'sd13))%(3'd7));
  localparam signed [3:0] p15 = {3{((2'd0)?(2'sd0):(3'sd0))}};
  localparam signed [4:0] p16 = ((~&(-3'sd2))?{1{(-2'sd1)}}:{4{(2'd1)}});
  localparam signed [5:0] p17 = ({2{(2'sd0)}}+(-(-5'sd3)));

  assign y0 = ($signed((((p14*a3)&(a2>=a4))))|$signed((((a3%b2)^(b5|p1)))));
  assign y1 = (({(a3^~b2)}^{3{b2}})|{4{{b5,a1}}});
  assign y2 = $unsigned({4{$signed($unsigned($unsigned($unsigned(p5))))}});
  assign y3 = (((p13&a4)?(a2===b5):{{b3}})<={(4'd6)});
  assign y4 = (&{1{($signed(((a3?a0:b4)?(b2>=b5):(-4'sd6))))}});
  assign y5 = (^((&({p1,b4}?(a1>p13):(~a0)))&((p4?p7:a1)?(|a1):{b5,p7,p9})));
  assign y6 = (5'd2 * (p12^~b2));
  assign y7 = (p1>a0);
  assign y8 = $unsigned((-(~|$unsigned(((4'd2 * (6'd2 * p2)))))));
  assign y9 = {1{{1{((a5)>>(b4===b1))}}}};
  assign y10 = (&p4);
  assign y11 = (!(&(~|(((a0===a3)>>>(&p16))<=((~|b1)>>>(p5-p14))))));
  assign y12 = {2{((b5+p4)+(p5>p9))}};
  assign y13 = (&((5'd9)|$unsigned((2'sd0))));
  assign y14 = (p4>b5);
  assign y15 = {(4'sd4),(2'd1),(5'd28)};
  assign y16 = ({1{{1{(((a4>=b1)||(b4&b4))==={4{b4}})}}}}||{4{{2{p5}}}});
  assign y17 = $unsigned((-$signed((~|(({b1,p16}==(b2>>p4))<={3{(b2-a5)}})))));
endmodule
