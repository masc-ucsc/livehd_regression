module expression_00582(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^(4'd2 * (4'd3)));
  localparam [4:0] p1 = {2{(((3'd3)<=(-4'sd7))===((5'd28)>(3'sd1)))}};
  localparam [5:0] p2 = ((2'd2)?(3'd4):(2'd2));
  localparam signed [3:0] p3 = ((~&{(~{2{{(4'sd1),(-3'sd2)}}})})>=(-{4{(4'd14)}}));
  localparam signed [4:0] p4 = ((((2'd2)?(4'd10):(3'd4))^~((2'sd0)?(4'd15):(2'sd0)))?(^((-3'sd3)<=(-5'sd3))):((4'd7)?(4'd9):(4'd6)));
  localparam signed [5:0] p5 = {((-5'sd7)?(3'd2):(4'd0)),{2{(5'sd8)}}};
  localparam [3:0] p6 = {(3'd6),{(5'd24)},((2'd0)?(5'd12):(5'd4))};
  localparam [4:0] p7 = {1{({1{((2'd0)!=(4'd1))}}<<<(((-5'sd3)|(5'd19))<((4'd14)<=(4'd4))))}};
  localparam [5:0] p8 = (-2'sd1);
  localparam signed [3:0] p9 = (&(~|((6'd2 * (4'd6))?(~^(-(2'sd0))):((3'sd3)+(2'd3)))));
  localparam signed [4:0] p10 = (3'd6);
  localparam signed [5:0] p11 = (((-5'sd11)&(5'd15))!==((-2'sd0)<<<(2'sd0)));
  localparam [3:0] p12 = (((4'sd2)&&(5'd14))?(2'sd0):((2'sd1)?(-5'sd8):(4'd14)));
  localparam [4:0] p13 = (~(|(~^(-(~|{2{(2'd2)}})))));
  localparam [5:0] p14 = (((3'd6)>=(+(3'sd1)))+(5'd31));
  localparam signed [3:0] p15 = (-5'sd5);
  localparam signed [4:0] p16 = ((3'sd2)>>>(|(4'sd4)));
  localparam signed [5:0] p17 = (~&(!(~^(({4{(-2'sd0)}}>=((2'd2)+(-4'sd2)))^~{1{(~&((4'd6)>=(4'sd2)))}}))));

  assign y0 = ({3{p12}}&&($signed($signed(p12))));
  assign y1 = (((5'd2 * p14)>>$unsigned((p8|p3)))<{((~|b5)),(p1|p10)});
  assign y2 = (5'sd2);
  assign y3 = (-3'sd3);
  assign y4 = ((a3!==a0)<{p4,p7});
  assign y5 = ({p6,a1,p2}||{p15,p15});
  assign y6 = (4'd2 * (4'd2 * b0));
  assign y7 = (a1===b0);
  assign y8 = $unsigned({2{{(!b0),{p3,a5}}}});
  assign y9 = {4{a1}};
  assign y10 = {2{(4'd9)}};
  assign y11 = (+($signed(((a3?p14:a3)>=(p6?p9:p2)))!=($unsigned(p17)^~(p1&&b2))));
  assign y12 = {1{((~(~^{2{(~&$unsigned((b0>b4)))}})))}};
  assign y13 = (((p0%b3)%p15)?((p14?b5:p4)>>>(a3?p1:p6)):((p10^a2)?(a5?a3:b0):(p2<p2)));
  assign y14 = ((+(b3>>a5))^((a4>a5)!==(a1?b0:b4)));
  assign y15 = (+(-4'sd3));
  assign y16 = (((b4>=a2)<{p15,a1})^{({a4}<=(a0<b0))});
  assign y17 = (^(-(~(-2'sd1))));
endmodule
