module expression_00112(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(^(4'd13)),((-5'sd1)+(2'd1)),(~(5'd16))};
  localparam [4:0] p1 = ((~(((3'd1)>>>(5'd0))<<{4{(5'd5)}}))?({4{(3'd3)}}?{3{(2'd1)}}:((3'sd1)>(4'd3))):(-{4{(2'd0)}}));
  localparam [5:0] p2 = ({1{{2{{4{(4'd7)}}}}}}<<<{1{(((5'd6)===(-2'sd0))==((3'sd2)^~(2'd0)))}});
  localparam signed [3:0] p3 = ((5'd31)<(2'sd0));
  localparam signed [4:0] p4 = (4'd2 * ((5'd1)?(5'd24):(4'd0)));
  localparam signed [5:0] p5 = (~(5'd30));
  localparam [3:0] p6 = {3{((5'd3)?(4'd11):(5'd29))}};
  localparam [4:0] p7 = ({(3'd7),(5'sd4)}?{(-5'sd9),(4'd7)}:((2'd2)?(4'd14):(-2'sd0)));
  localparam [5:0] p8 = {3{((-2'sd1)?(5'd2):(2'd2))}};
  localparam signed [3:0] p9 = {1{{4{(2'd1)}}}};
  localparam signed [4:0] p10 = ((~|{(-{(2'd2),(2'd2)}),((4'd6)!=(5'sd9))})||({{3{(-2'sd0)}}}==((2'd2)|(-2'sd1))));
  localparam signed [5:0] p11 = {4{{(3'd4),(5'sd1),(-2'sd1)}}};
  localparam [3:0] p12 = (4'sd4);
  localparam [4:0] p13 = ((&((4'd3)?(2'sd0):(2'd2)))&({3{(5'sd14)}}^(4'd2 * (4'd9))));
  localparam [5:0] p14 = {3{(|(5'sd2))}};
  localparam signed [3:0] p15 = {2{(-4'sd5)}};
  localparam signed [4:0] p16 = (((((2'd3)===(5'd13))>>>((3'd7)+(5'd11)))>(((4'd3)/(5'd17))>>>((2'd1)<<(-5'sd8))))!=((((5'sd15)<=(-3'sd3))/(-2'sd0))>>(5'd2 * ((3'd1)===(3'd5)))));
  localparam signed [5:0] p17 = (+{(-(2'sd0))});

  assign y0 = (5'sd9);
  assign y1 = {4{p17}};
  assign y2 = {1{{3{({2{a3}}<<(p5-b0))}}}};
  assign y3 = {p15,p6,p12};
  assign y4 = {b5,b1,b2};
  assign y5 = {1{{(3'd3),{3{{3{p16}}}},((5'd19)<<{p10,p13})}}};
  assign y6 = (~^(5'sd2));
  assign y7 = (2'd1);
  assign y8 = (({((a5!==a2)?{p5,p13,p10}:(~|a0)),(|(a1?p1:p2)),(-(~^((p2?a2:b4))))}));
  assign y9 = (2'd2);
  assign y10 = $unsigned({({$unsigned(a4),(-4'sd0)}^~$signed((2'd1)))});
  assign y11 = (((a0?a1:p4)?(b5?p13:p8):(b5?p15:p12))?{{(p13?p0:p6),(p16?p9:a4)}}:{(a1?p14:p7),{p8,p10,p6}});
  assign y12 = (6'd2 * (a0>=b0));
  assign y13 = {2{(p0?p11:a1)}};
  assign y14 = (p14>>p5);
  assign y15 = $unsigned((&(p1)));
  assign y16 = ({(p12<<p10),(2'sd1),(!(|p10))}>>(-3'sd2));
  assign y17 = ((2'sd1)?({p13}?{p14,p4,p14}:(|p1)):((p5?p11:p3)?(&p0):(p0?p0:p15)));
endmodule
