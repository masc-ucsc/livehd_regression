module expression_00669(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd0)*(-4'sd2))&((2'd0)||(2'd0)))|(((5'd2)<<(2'd1))?((5'sd3)!==(3'sd2)):((-3'sd1)>(5'd12))));
  localparam [4:0] p1 = {3{(((4'sd2)&&(-5'sd11))<<<((2'sd1)<(-2'sd1)))}};
  localparam [5:0] p2 = ({{1{(2'd0)}},((-3'sd3)>>(-3'sd3))}==(((4'd12)===(5'sd7))>(|(5'sd4))));
  localparam signed [3:0] p3 = (4'sd6);
  localparam signed [4:0] p4 = (((-5'sd2)<<<(2'd2))?(4'sd6):{1{((5'sd12)?(5'd27):(-3'sd3))}});
  localparam signed [5:0] p5 = (^(~&{1{(((4'sd2)?(5'd14):(5'sd12))===(~&(3'sd0)))}}));
  localparam [3:0] p6 = ((((5'd1)|(-5'sd5))&&((4'd7)&(4'd7)))?(((5'd1)<(3'd0))^{3{(5'd16)}}):{3{((5'sd10)<(2'd0))}});
  localparam [4:0] p7 = ((-3'sd0)*(5'd25));
  localparam [5:0] p8 = (|(~(3'd4)));
  localparam signed [3:0] p9 = (3'sd2);
  localparam signed [4:0] p10 = ((((2'sd0)>>(5'd16))<<((4'd13)>(4'sd1)))||({(-4'sd0),(-4'sd1),(4'd14)}^((4'd15)&(3'd1))));
  localparam signed [5:0] p11 = ((2'd1)>=((3'sd1)===(-2'sd0)));
  localparam [3:0] p12 = {1{{1{(+((~&(+(-5'sd3)))?{4{(2'd1)}}:{(3'sd0),(5'sd12)}))}}}};
  localparam [4:0] p13 = ((-4'sd3)==(5'd10));
  localparam [5:0] p14 = ((3'sd1)!=(3'd0));
  localparam signed [3:0] p15 = {(^(3'd2))};
  localparam signed [4:0] p16 = (3'd2);
  localparam signed [5:0] p17 = (({3{(3'd6)}}<<(5'd2 * (3'd7)))<<{3{{1{(-3'sd2)}}}});

  assign y0 = ({2{(~&{3{{3{p13}}}})}});
  assign y1 = {{p14,a2,p17},(b0?p12:a2)};
  assign y2 = {4{({p16,b4}+{b0,p13,b1})}};
  assign y3 = (($signed((-p10))^~(b3?a3:a2))!=({2{b5}}+$unsigned((a2?p8:b4))));
  assign y4 = (({1{$signed(($signed((b5?b3:b4))))}})?({4{a5}}?$signed(a4):(b4?a0:p4)):{4{(b5)}});
  assign y5 = (5'd29);
  assign y6 = (~&(~^(a4)));
  assign y7 = (2'd1);
  assign y8 = {(~&({({b2,b1,p12}|(p1+p4))}&&(!(!{(2'd0)}))))};
  assign y9 = {{(-5'sd11)}};
  assign y10 = (!{((-(~^(~|((p15|p10)||(p0+p11)))))&((&(p11<=p5))<<(-(+(p7<p11)))))});
  assign y11 = ((~^a2)>>$unsigned(p0));
  assign y12 = (a3?a1:b0);
  assign y13 = (((a4<b0)<<<(b2^a2))===(|((b1!==b0)<(b0===b1))));
  assign y14 = ((a5^~p0)^~(3'd2));
  assign y15 = {4{{4{p9}}}};
  assign y16 = (~(((p12^~p15)?{4{p4}}:{b1})?{(~^b3),{b1,a4,p16},(p10>>b4)}:(-(p0?p2:p7))));
  assign y17 = ((p1<p7)<=$unsigned($signed(p0)));
endmodule
