module expression_00847(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(|((|(!((!(4'd3))*((-4'sd7)|(4'sd3)))))||(+(^(+(((-5'sd8)+(3'sd2))>((-3'sd1)/(-2'sd0)))))))));
  localparam [4:0] p1 = ((-4'sd7)?(-2'sd1):(2'd2));
  localparam [5:0] p2 = {(({{(-3'sd0),(-4'sd1)}}>((-2'sd1)?(-2'sd0):(5'd31)))&{((5'd28)||(2'd3)),((2'sd1)?(-4'sd7):(5'sd5))})};
  localparam signed [3:0] p3 = (4'd6);
  localparam signed [4:0] p4 = ((((2'd2)?(2'd2):(3'd2))?((-3'sd0)||(-5'sd11)):(4'd2 * (4'd5)))^(((5'd4)?(4'd4):(3'd0))|((5'd27)?(2'd1):(2'd3))));
  localparam signed [5:0] p5 = ({(&(2'd0)),{3{(-5'sd9)}},((5'sd8)<=(-4'sd4))}^{(~&{(|{4{(3'd4)}})})});
  localparam [3:0] p6 = (3'sd2);
  localparam [4:0] p7 = (({(3'd1),(3'sd1),(-2'sd1)}!={(5'd17)})?{3{(~(4'd10))}}:{2{(+(5'd6))}});
  localparam [5:0] p8 = (~^(~&{{{(2'd3),(3'd7)},(-(-2'sd1)),{(3'd3),(5'd14),(5'd3)}}}));
  localparam signed [3:0] p9 = (((2'sd1)&&(2'sd0))?(~&(5'd8)):((4'd12)!==(2'd0)));
  localparam signed [4:0] p10 = (^((-((^(-4'sd5))<=((5'd5)?(4'd11):(3'd6))))>>>(!(!(((4'sd1)<<<(3'sd3))&(|(4'd6)))))));
  localparam signed [5:0] p11 = {(5'sd10)};
  localparam [3:0] p12 = ((-4'sd2)+((-2'sd0)/(2'sd1)));
  localparam [4:0] p13 = {(-3'sd1),(-2'sd1)};
  localparam [5:0] p14 = (~(~^(&(4'd1))));
  localparam signed [3:0] p15 = (((3'd0)?(3'sd1):(-3'sd3))>(-4'sd5));
  localparam signed [4:0] p16 = {{(2'd2),{(-4'sd5)}},(~&{1{{(2'd1),(5'd27)}}}),(-2'sd1)};
  localparam signed [5:0] p17 = (~^(5'd5));

  assign y0 = (|({4{(p13&&p1)}}||(((~|p0)<=(!p2))||{1{{2{a3}}}})));
  assign y1 = {{(+(p3<p8))},{2{{p0,p16,p12}}},(|(p1^~p5))};
  assign y2 = (+(~|(-($unsigned((^(+({p12}&&(~^p9)))))<<(-5'sd14)))));
  assign y3 = ((a3?b3:b5)!==(a2-b4));
  assign y4 = {1{(({3{b5}}!==(b0<<<b2))<<<(p11?p13:p11))}};
  assign y5 = {3{((p16)-{p12,p6,p7})}};
  assign y6 = {2{((b0)||(~|a3))}};
  assign y7 = (+(+((~|(b3>>>b0))>(&(&(+b4))))));
  assign y8 = ($unsigned(({(p16?a5:p6),(p14?p5:b3)}?(p13?a4:b3):$unsigned((b0?b4:a2)))));
  assign y9 = {2{(b3-b0)}};
  assign y10 = (3'sd0);
  assign y11 = ((~&(((p7||p3))<(p5<<<p11)))^~(((~p16))|(3'sd2)));
  assign y12 = (b4?a1:p7);
  assign y13 = (~&((3'd4)!=$unsigned(($signed(({2{p3}}=={2{b3}}))))));
  assign y14 = (~|{p2});
  assign y15 = ((((a0^a1)<={3{a2}})===(~^(b5|b4)))-{1{{3{(a5<<<a5)}}}});
  assign y16 = (p3?p16:p13);
  assign y17 = (~(5'd27));
endmodule
