module expression_00270(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd2)?{4{(3'd6)}}:(5'sd5));
  localparam [4:0] p1 = (~|(2'sd0));
  localparam [5:0] p2 = (((2'd1)<(4'd15))==(~((-3'sd0)>=(3'd0))));
  localparam signed [3:0] p3 = (&(~(+((&(4'd9))>>{4{(2'd1)}}))));
  localparam signed [4:0] p4 = {{3{{(-4'sd5)}}},(!{3{(3'sd2)}})};
  localparam signed [5:0] p5 = {{(-5'sd8),(5'd29),(2'd3)}};
  localparam [3:0] p6 = {2{(2'sd1)}};
  localparam [4:0] p7 = ((^(3'sd3))^(|(3'd7)));
  localparam [5:0] p8 = (2'd0);
  localparam signed [3:0] p9 = (({2{(3'sd2)}}?(-(2'sd1)):(~(5'd29)))?({2{(3'd1)}}?((5'd18)||(4'd11)):(~&(-3'sd0))):((~|(3'd2))?(~^(-2'sd1)):(~&(3'sd2))));
  localparam signed [4:0] p10 = {4{{3{(5'sd13)}}}};
  localparam signed [5:0] p11 = (-3'sd3);
  localparam [3:0] p12 = {4{((-5'sd4)^~(4'd9))}};
  localparam [4:0] p13 = {{{{(2'sd0),(2'd1),(5'd13)},(|(-5'sd0)),((3'sd1)?(3'd3):(-2'sd0))}},(^{(-(-3'sd0)),((-4'sd4)?(2'd0):(5'd14)),(~(3'd5))})};
  localparam [5:0] p14 = ((5'd22)?((-5'sd5)?((-4'sd3)?(3'd6):(4'd1)):(5'sd15)):(((2'd3)^(4'sd3))==(5'sd6)));
  localparam signed [3:0] p15 = ({(5'd25),(3'd7)}?(|(-4'sd6)):((2'd2)?(-4'sd7):(-2'sd1)));
  localparam signed [4:0] p16 = (({4{(5'd17)}}-((3'd2)^~(2'd0)))&((5'd2 * (3'd6))>>>{3{(2'd1)}}));
  localparam signed [5:0] p17 = (((-2'sd0)<<<(3'sd3))?((2'd2)?(4'd15):(5'd31)):((-2'sd1)?(-3'sd2):(2'd0)));

  assign y0 = (((-5'sd9)<(b2&&a2))!==(2'sd0));
  assign y1 = (b3?p14:p1);
  assign y2 = (-3'sd0);
  assign y3 = $unsigned((-3'sd2));
  assign y4 = ((+{2{((~^{1{{2{p12}}}})>>>{3{p17}})}}));
  assign y5 = (-2'sd1);
  assign y6 = ($signed((&p2))^(a3<<<p5));
  assign y7 = ({3{b2}}===(&{b1,a1,b3}));
  assign y8 = (~^(|(((^$signed((2'd1))))?(^(|(4'sd5))):((3'sd3)?$unsigned(p0):(p17?p17:p0)))));
  assign y9 = (5'd9);
  assign y10 = {1{(3'd4)}};
  assign y11 = ({((($unsigned(p3))<<<(5'sd4))<<<($unsigned({{b0,b5},$unsigned(b0)})))});
  assign y12 = (((4'sd1)>=(-((p0+a0)|(p9^b0))))!=(6'd2 * (2'd0)));
  assign y13 = ((a3==b4)&(b2?a0:a5));
  assign y14 = (p10|p7);
  assign y15 = (b3?p10:p10);
  assign y16 = {$unsigned({p5,p9}),{(-4'sd6)},$signed({p9,b2,p4})};
  assign y17 = ((p3?b5:p12)?(p11?p8:a3):(p8<<p11));
endmodule
