module expression_00358(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({2{{1{((4'd3)?(-4'sd3):(3'd2))}}}}&((-(3'd0))?{2{(2'd3)}}:{3{(-4'sd1)}}));
  localparam [4:0] p1 = (~^(!(-((-5'sd10)?{2{(5'sd2)}}:(~|(2'd1))))));
  localparam [5:0] p2 = (2'd1);
  localparam signed [3:0] p3 = (((5'd3)&(2'sd0))<(!((2'sd1)>=(-3'sd1))));
  localparam signed [4:0] p4 = (3'd2);
  localparam signed [5:0] p5 = (3'sd0);
  localparam [3:0] p6 = {{1{(-5'sd2)}},(2'd1)};
  localparam [4:0] p7 = {3{(!(5'sd0))}};
  localparam [5:0] p8 = (({((5'sd7)!==(2'sd0)),((-3'sd0)<<<(2'sd0))}&(((3'sd3)===(4'sd3))>=((-5'sd1)>=(2'd2))))<<({(2'd3),(2'sd0),(-4'sd7)}==(((-5'sd6)&(-5'sd8))=={(2'sd1),(2'd2)})));
  localparam signed [3:0] p9 = (((-2'sd1)?(2'sd1):(5'd10))?(5'sd1):(-2'sd0));
  localparam signed [4:0] p10 = ((6'd2 * (3'd0))?((5'sd7)?(2'd2):(3'd6)):(2'sd1));
  localparam signed [5:0] p11 = (&(~&(~|(5'sd12))));
  localparam [3:0] p12 = {4{((-2'sd1)+(3'd7))}};
  localparam [4:0] p13 = ({2{(~(3'sd3))}}+((4'd2 * (5'd4))!==((2'd1)<=(4'd3))));
  localparam [5:0] p14 = ((((4'sd4)^~(2'd2))?(~^((4'sd5)?(-4'sd1):(2'sd0))):((3'sd2)?(-5'sd2):(-4'sd6)))^(6'd2 * ((3'd0)^(4'd5))));
  localparam signed [3:0] p15 = ((((4'd7)<<<(2'd2))!=(~|(-2'sd0)))?(((3'd6)>=(-2'sd1))||((-4'sd2)===(-4'sd5))):((~^(-5'sd14))==((5'sd10)?(3'd6):(4'd1))));
  localparam signed [4:0] p16 = ((-3'sd1)-(-3'sd0));
  localparam signed [5:0] p17 = ({2{((2'sd0)?(4'sd2):(2'd1))}}<=((-3'sd0)?(4'd15):(5'd1)));

  assign y0 = (($signed(((b5)===(a3&&a0)))<<((b0!==b1)?(p1?a0:b5):(b2?a3:a3)))<<<((b1?a0:p0)?$unsigned((b0===b4)):$signed($unsigned(a0))));
  assign y1 = (a4?b4:b2);
  assign y2 = (&(($signed((((3'd7)>>(p16||b4))+(2'd0))))<(5'sd13)));
  assign y3 = (((p1?p12:p2))?(a2?b0:a5):(p8?b4:p9));
  assign y4 = (b5+p6);
  assign y5 = (3'd4);
  assign y6 = ((~|(-((b2?a4:b4)===(!b2))))?((~&(|p11))|(&(p6?b1:p16))):(~((|(!p17))!=(~&(~a4)))));
  assign y7 = (4'd13);
  assign y8 = (+(5'd2 * {(p7?p6:p8)}));
  assign y9 = {4{(&a0)}};
  assign y10 = ((~|((b1?a0:p15)^~((b2?b1:a2)+(b5?a5:p12))))&(|(~^(~^((^(b0>b2))!==(b4?a4:a1))))));
  assign y11 = (-4'sd6);
  assign y12 = {4{{3{a0}}}};
  assign y13 = (~{1{(+(|$signed($unsigned({2{{3{b2}}}}))))}});
  assign y14 = (+((~^{{(&b2)},(^(a0&&b0)),(~|(-4'sd0))})>((6'd2 * {a2})<=(|(|(p7+b0))))));
  assign y15 = (|({3{(3'd5)}}||{3{(b3===b0)}}));
  assign y16 = (-{({b1,a1,p7}>>(p16^p17)),{1{(3'sd2)}},(|(2'sd0))});
  assign y17 = (4'd8);
endmodule
