module expression_00556(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-3'sd0)?(2'd2):(2'd0));
  localparam [4:0] p1 = {1{({2{{4{(-5'sd3)}}}}>=({3{(3'd1)}}>=((4'd3)?(5'd7):(4'd2))))}};
  localparam [5:0] p2 = ((3'sd1)?(-5'sd5):(-4'sd4));
  localparam signed [3:0] p3 = ((|(~(3'sd3)))?((4'sd6)>>(2'sd1)):(^((2'd1)?(4'd10):(2'd2))));
  localparam signed [4:0] p4 = ({1{((4'sd4)&&(4'd7))}}+((4'sd3)!=(2'sd1)));
  localparam signed [5:0] p5 = {(-4'sd2),{{(5'd6)}},(3'd2)};
  localparam [3:0] p6 = ((4'sd4)!=((3'sd2)>=(3'sd0)));
  localparam [4:0] p7 = (((3'd2)==(3'd3))+((2'd0)>(2'sd1)));
  localparam [5:0] p8 = (-(&((+((~&(2'sd0))!==((2'd1)+(5'd30))))!=(!(|(-((5'd21)!=(5'sd0))))))));
  localparam signed [3:0] p9 = {((|(~(4'd8)))==={4{(3'sd1)}}),(~&((4'd8)==={3{(-5'sd8)}}))};
  localparam signed [4:0] p10 = (((|(-5'sd2))?(~(-4'sd3)):((-2'sd1)?(5'sd13):(-4'sd7)))?(~|{(5'd13),(4'sd2),(-4'sd2)}):(((5'd14)?(4'sd0):(3'd0))?{(5'sd0),(3'd7)}:(&(3'd7))));
  localparam signed [5:0] p11 = ((((4'd1)?(5'd13):(4'd7))?(&(3'd3)):(-4'sd7))>=(5'd18));
  localparam [3:0] p12 = {1{((5'd29)=={3{(-4'sd4)}})}};
  localparam [4:0] p13 = (3'd7);
  localparam [5:0] p14 = ((-4'sd3)>>(-3'sd1));
  localparam signed [3:0] p15 = (((3'sd3)?(2'sd1):(-2'sd1))?{(-3'sd3),(2'sd0)}:{(3'sd3)});
  localparam signed [4:0] p16 = (((2'd2)?(-5'sd10):(4'd4))<<<(((3'sd1)<=(2'd0))^((4'd4)>>(3'd0))));
  localparam signed [5:0] p17 = (((-4'sd2)<(-2'sd1))*(-((3'd3)||(3'd7))));

  assign y0 = (-(-2'sd1));
  assign y1 = ((~&(~(p2?p9:p4)))?(!(a2?p8:p2)):(b5?p13:p13));
  assign y2 = (4'sd7);
  assign y3 = ((~|(-3'sd3))/a0);
  assign y4 = {(4'sd3),(&{3{p11}})};
  assign y5 = {{{a0},{b3,p13},{p17,p12,b3}},({{p10,p0}}&(p13>>>p10)),({a1,p13,b4}<={b1,a3,p1})};
  assign y6 = $signed($unsigned($signed($unsigned(p1))));
  assign y7 = (~^{b3,a3,b5});
  assign y8 = ((p9!=a0)?(a4^p1):(p1?p11:p6));
  assign y9 = (!((a3+p14)+{2{a1}}));
  assign y10 = {4{(~&(!p14))}};
  assign y11 = ((~|(-(p13?p9:p16)))?((p8?p9:p1)?(p6?p3:p10):(-p16)):((p14<<p1)?(p12==p9):(5'd2 * p13)));
  assign y12 = {(((p9?p1:p7)?(p13>=p10):(p17?p7:p4))==(((p12^p3)&&(p6^p2))>>{p5,p0,p0}))};
  assign y13 = (^((~(~&p7))&&(~&(a3<<p8))));
  assign y14 = ((((b4%a3)%a0)==(~(~&(a2===b3))))>>(((-a2)^~(a0&a1))|(&(p1<<<a1))));
  assign y15 = (((~({a3}^~(~b5)))!==((a5|b4)-(b4^~a2)))|((^(4'd2 * {p12,p12,p13}))!=({2{a5}}&(p9<<a0))));
  assign y16 = {2{({1{(~|p12)}}|{2{p11}})}};
  assign y17 = (-(({2{b0}}>={(a0?b5:b3)})<{2{{3{a3}}}}));
endmodule
