module expression_00121(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd2)||(3'sd3));
  localparam [4:0] p1 = (4'd2);
  localparam [5:0] p2 = (((4'd2 * (4'd15))>=(5'd2 * (2'd1)))>>(((4'd5)?(-5'sd8):(-5'sd13))?((5'd24)?(-4'sd5):(-2'sd1)):((5'd0)?(-3'sd0):(3'd4))));
  localparam signed [3:0] p3 = (~|((-3'sd2)?(5'd15):(5'd11)));
  localparam signed [4:0] p4 = {(3'd0)};
  localparam signed [5:0] p5 = {4{(((4'd11)!=(3'd2))-((3'd7)>=(5'd3)))}};
  localparam [3:0] p6 = ((5'd31)&(-3'sd0));
  localparam [4:0] p7 = ({2{(4'd7)}}?(|(~^(3'd3))):(~(|(-3'sd0))));
  localparam [5:0] p8 = ((2'sd0)?(5'd18):(-4'sd5));
  localparam signed [3:0] p9 = (-3'sd1);
  localparam signed [4:0] p10 = {3{((-3'sd0)!==(3'd3))}};
  localparam signed [5:0] p11 = {(~|(~^(4'sd4))),{{(5'd6)}},((3'd7)^(-4'sd5))};
  localparam [3:0] p12 = (~&(~(^(2'sd1))));
  localparam [4:0] p13 = (~&((~^((-5'sd7)?(-3'sd1):(2'd1)))?(!((5'd1)&&(2'd1))):((|(2'd0))|((-2'sd0)-(-4'sd7)))));
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = (-5'sd11);
  localparam signed [4:0] p16 = ((((5'd27)-(3'd6))?((2'd2)?(-3'sd0):(-2'sd0)):((-5'sd5)!=(3'd7)))+(((3'd2)?(2'd3):(5'sd9))?{2{(4'sd5)}}:((-4'sd1)?(2'd1):(4'd1))));
  localparam signed [5:0] p17 = ((((2'd2)>=(4'd4))===((-4'sd4)&(4'd9)))<<<{((-2'sd1)<<<(-2'sd1)),((5'd20)<(2'sd0)),((-3'sd2)^~(3'd2))});

  assign y0 = ({4{a3}}?{2{(5'd2 * p0)}}:{{1{(p2?b4:p15)}}});
  assign y1 = $signed(p11);
  assign y2 = ((a1&p1)?{p2,p4,b0}:(|a0));
  assign y3 = (^$signed(((&(({3{b0}}<={2{b0}}))))));
  assign y4 = (b5?p2:b3);
  assign y5 = (~|$unsigned(((~|b4)||$unsigned(p15))));
  assign y6 = ((4'd8)?((-b4)?(p11?a0:a3):(a1^~p10)):((-(3'd6))>(3'd0)));
  assign y7 = (~|(-{1{(~|(-5'sd0))}}));
  assign y8 = (|(~&(~(+{(-({((p3?p3:p10)<=(~&(a5!==a4)))}<<((a5||b4)?(b3==b3):(p7?b0:a1))))}))));
  assign y9 = {$signed((~p14)),(a5?p1:b2)};
  assign y10 = ((3'd6)!==(2'sd1));
  assign y11 = {$signed((3'sd2))};
  assign y12 = (2'sd0);
  assign y13 = {3{((p15?p5:p16)?(a5&&a5):(a4<<a0))}};
  assign y14 = ((~|({3{p14}}>>{4{p8}}))>{2{((p4+p14)-(p9>>p9))}});
  assign y15 = (|((+p13)&$signed(b2)));
  assign y16 = (5'd30);
  assign y17 = ({{{p2},(p16?p15:p16),(p1?p0:p8)}}?{({p14,p13,p0}?{p12}:(p13?p7:p5))}:{{p10,p10},(p7?p9:p13)});
endmodule
