module expression_00664(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^{((2'd2)>>((5'd30)^(4'd14)))});
  localparam [4:0] p1 = ((4'd0)?(5'd17):(4'd2));
  localparam [5:0] p2 = (((2'd0)<=(3'd6))||((2'd2)>>>(2'sd0)));
  localparam signed [3:0] p3 = {{1{{2{(5'd19)}}}}};
  localparam signed [4:0] p4 = ((((2'sd1)?(3'd4):(-3'sd3))||((-4'sd2)<<<(-5'sd13)))?(((5'sd1)<=(3'sd0))===((3'd0)?(-5'sd6):(3'd7))):(((-4'sd0)&(-3'sd1))^((3'd6)?(-4'sd3):(2'sd1))));
  localparam signed [5:0] p5 = (|(&(!(-(&(~|{1{{2{{2{(2'd2)}}}}}}))))));
  localparam [3:0] p6 = (((-2'sd1)|(3'd7))?{(3'd5),(2'd2),(3'd6)}:((5'sd15)!=(2'd0)));
  localparam [4:0] p7 = (|((&{2{(4'sd0)}})>{(5'd4),(5'd13)}));
  localparam [5:0] p8 = {{3{(4'd11)}},(((4'd7)<<(-4'sd0))==={(5'sd15),(2'd3),(2'd1)})};
  localparam signed [3:0] p9 = ((4'sd2)!==({2{(2'd3)}}?(~&(2'd1)):(&(5'd25))));
  localparam signed [4:0] p10 = ({{(5'd21)},(~^(3'd7)),(!(5'd19))}?{(~|(~^((-4'sd0)!=(-5'sd7))))}:(|((~^(5'd29))!=(!(2'd1)))));
  localparam signed [5:0] p11 = (-3'sd1);
  localparam [3:0] p12 = (((-3'sd1)?(-2'sd0):(-5'sd12))?(2'd1):((5'd24)<<<(3'd1)));
  localparam [4:0] p13 = (2'd2);
  localparam [5:0] p14 = ({4{(-3'sd0)}}+{(4'sd5),(2'd1)});
  localparam signed [3:0] p15 = (&(^(((~&(4'd15))>>(-(5'd16)))?{{((5'd0)|(2'd3))}}:(!((5'sd3)&&(5'd17))))));
  localparam signed [4:0] p16 = ((2'd3)/(-2'sd0));
  localparam signed [5:0] p17 = (!(({(5'd3)}>{(3'd4)})-{((4'd5)^(-3'sd0)),((5'sd1)&&(5'sd10)),{(4'd10),(2'sd0),(4'd0)}}));

  assign y0 = ((b1?a5:a1)?(b1?b5:b5):(a1<<b1));
  assign y1 = (!{{1{(~^((!{2{b1}})&{4{a5}}))}}});
  assign y2 = (5'd5);
  assign y3 = (((p9?b4:p6)%p1)^($unsigned((p1?p15:p14))&(p15?p8:p5)));
  assign y4 = (2'sd0);
  assign y5 = ((~&(&(~&(p4?b1:b4))))>>>(-(~|{1{(b5&&b2)}})));
  assign y6 = ((3'd7)?(4'd4):(4'sd1));
  assign y7 = ((4'd15)<<(4'd2 * (b2|p7)));
  assign y8 = {$unsigned((|(&({(p17^~a1),(|p8)}))))};
  assign y9 = $unsigned((((p16==b3)||(b4?a5:a3))?(+((+b5)<<(-p17))):((p17?p9:p10)<<(~|p7))));
  assign y10 = (^$signed((~(({1{p3}}&{1{a0}})|(-{3{p16}})))));
  assign y11 = (((|a3)?(b3?a3:b4):(~|a5))?((~a4)?$unsigned(a3):(^b2)):((|p7)?(~b2):(a0?p8:b3)));
  assign y12 = (5'sd3);
  assign y13 = (-2'sd1);
  assign y14 = (((a1===b3)?(~^a3):(a3>>>a5))!==((3'd3)?(5'd17):(-4'sd7)));
  assign y15 = ((-(~^(b4*a3)))||(|(&(^(!a2)))));
  assign y16 = {(+p0),{p17},(~&p10)};
  assign y17 = ({4{(a3!==a5)}}-{1{{3{{3{a0}}}}}});
endmodule
