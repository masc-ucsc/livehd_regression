module expression_00097(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(~&((3'd5)?(2'd2):(-5'sd11))),((2'd3)?(2'sd0):(5'd10)),(~^(|(~|(-4'sd2))))};
  localparam [4:0] p1 = ((!(-(-5'sd5)))<{3{(4'sd3)}});
  localparam [5:0] p2 = ({3{(3'd2)}}<<((5'sd4)+(3'd2)));
  localparam signed [3:0] p3 = (({3{(-2'sd0)}}>>>(6'd2 * (5'd31)))>=((^(5'd9))>((3'sd2)?(5'd17):(2'd2))));
  localparam signed [4:0] p4 = {3{(3'd1)}};
  localparam signed [5:0] p5 = {4{{(4'd4),(4'd11)}}};
  localparam [3:0] p6 = ((4'd14)?(3'd5):(5'd0));
  localparam [4:0] p7 = (4'd2 * (5'd19));
  localparam [5:0] p8 = (((5'd2 * (2'd3))!=((4'd1)&&(5'd22)))^(~|(-((4'sd3)==(-4'sd5)))));
  localparam signed [3:0] p9 = (-{((2'd2)?(3'd7):(4'd11)),((4'd5)?(-2'sd0):(-5'sd9))});
  localparam signed [4:0] p10 = (((+((4'sd0)+(3'sd0)))&&((5'd26)==(4'd15)))!==(!(((-4'sd1)!=(5'sd9))>>((3'd6)===(5'sd9)))));
  localparam signed [5:0] p11 = ((((-4'sd2)*(-2'sd1))%(4'd0))?(((4'd1)?(-2'sd0):(2'd0))?(~|(3'd2)):(~^(3'd6))):((~|((4'sd0)<<<(5'd22)))%(4'd12)));
  localparam [3:0] p12 = (3'd1);
  localparam [4:0] p13 = (~|(~|(((-5'sd10)===(5'd6))+(|(|(5'd2))))));
  localparam [5:0] p14 = ((~^((2'd0)?(3'd3):(4'd2)))>>>(~(^((3'd5)^~(3'd3)))));
  localparam signed [3:0] p15 = {4{(2'd0)}};
  localparam signed [4:0] p16 = (((4'sd7)||(-2'sd0))<=((3'sd2)?(3'd5):(-3'sd3)));
  localparam signed [5:0] p17 = (5'd10);

  assign y0 = {(a2?b1:a1),{{3{b2}}},(~|{4{b1}})};
  assign y1 = ((p12?p3:a4)>>{2{(p14<b3)}});
  assign y2 = ($signed({$unsigned(p4),(p16||p17)})-(5'sd13));
  assign y3 = (4'd2 * (6'd2 * b0));
  assign y4 = {((b4?p13:b4)?{p1,a0,b3}:{a1,a2}),((-{4{a5}})?{4{b1}}:{a3,a1,a2})};
  assign y5 = {4{(a5?a1:b5)}};
  assign y6 = (5'sd13);
  assign y7 = ((((^$signed(b3))&&(~{3{a1}}))^~(-{2{{3{p10}}}})));
  assign y8 = {{(b2|a3),(p0)},$signed(((4'd5)|(4'd8))),{{a2,a5,b0}}};
  assign y9 = (((p16?p13:a5)?(~&p10):(4'd8))?(6'd2 * (-(~|a1))):((|p9)?(p14*p10):(3'd4)));
  assign y10 = {2{(b5!=a5)}};
  assign y11 = (4'd5);
  assign y12 = (+(a3<<<p7));
  assign y13 = ({4{b5}}^{{a5,a4,p16}});
  assign y14 = $signed(({1{{1{(2'd1)}}}}));
  assign y15 = $unsigned($signed((($unsigned(($unsigned(p17)))))));
  assign y16 = $unsigned(({2{$signed((a0>=p16))}}^{4{(p4==p9)}}));
  assign y17 = ({4{(p8==p1)}}<(^((-2'sd0)!=((p13||p8)^{2{b5}}))));
endmodule
