module expression_00562(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(~|(-(((4'sd1)?(5'sd1):(4'd8))?((3'd6)?(4'd10):(2'sd1)):((5'sd10)?(-4'sd6):(-2'sd1))))));
  localparam [4:0] p1 = (~&(~(^((-4'sd4)>>(-3'sd1)))));
  localparam [5:0] p2 = (-(3'd1));
  localparam signed [3:0] p3 = (((3'd4)?(4'd15):(4'sd5))*((3'd7)-(2'd1)));
  localparam signed [4:0] p4 = ((~&((-((2'd0)?(3'sd3):(5'd19)))+(+((3'sd2)===(-2'sd0)))))>=(((-4'sd0)<=(-5'sd1))^(+((-4'sd4)&&(-5'sd9)))));
  localparam signed [5:0] p5 = {{((3'd3)?(2'd2):(-3'sd2))},{((4'sd7)===(5'd31))},((5'd14)>(3'd0))};
  localparam [3:0] p6 = {3{(-3'sd2)}};
  localparam [4:0] p7 = ({{(-2'sd0),(4'd9),(3'd2)},{(2'd1),(-5'sd7),(-3'sd2)}}?((-3'sd0)?(5'd28):(5'd24)):((4'd3)?(5'sd3):(3'd6)));
  localparam [5:0] p8 = (({(3'd5),(5'd18)}&(~|(-4'sd5)))?(&(~|((5'd31)>>>(2'd2)))):(((4'd4)?(3'sd3):(2'd0))<=((2'sd1)!==(4'sd0))));
  localparam signed [3:0] p9 = {((4'd10)!=(4'sd5)),{3{(2'sd0)}},{2{(2'd1)}}};
  localparam signed [4:0] p10 = (-{3{{2{{(4'd0)}}}}});
  localparam signed [5:0] p11 = (&(~&{{(2'd2),(5'sd11),(4'd8)}}));
  localparam [3:0] p12 = {(6'd2 * {(3'd7),(5'd12)})};
  localparam [4:0] p13 = (2'sd0);
  localparam [5:0] p14 = {1{(3'sd2)}};
  localparam signed [3:0] p15 = (!((5'd30)==((4'd7)<(~&((4'sd7)^~(3'sd3))))));
  localparam signed [4:0] p16 = ((-5'sd9)>>(-2'sd1));
  localparam signed [5:0] p17 = (~^((((5'sd9)>>>(2'sd1))==((-5'sd15)==(5'sd5)))<<(-((+(-5'sd4))?((3'd1)&(3'd6)):((4'd14)^(-4'sd3))))));

  assign y0 = ({1{((-a1)?{4{b3}}:(p6?p3:p4))}}?((a4)?(a3|p0):(p6?p2:a2)):$unsigned(((p9?a3:a5)?(b4|b3):(a4|p4))));
  assign y1 = (-3'sd1);
  assign y2 = {3{b3}};
  assign y3 = {4{(a0||p4)}};
  assign y4 = {(~(p10?p3:p5))};
  assign y5 = {4{a2}};
  assign y6 = ({b5,a2}===(b5^a0));
  assign y7 = (((p14+b3)^~$signed((a4)))?((a1?p7:a2)/a1):(~^((~|(b4|p15))!=$signed((~|a5)))));
  assign y8 = (4'd9);
  assign y9 = $signed($signed((a3?a2:a0)));
  assign y10 = ((p11?p11:p5)?{p3,p17,p12}:{4{p2}});
  assign y11 = ($unsigned(((|p15)||(p13<=p5)))&(5'sd2));
  assign y12 = ({(a0-b0),(~^(~&a5))}!=(~&(3'd2)));
  assign y13 = {{(2'd3),$signed((4'sd6))},(((p0?p7:b5))-(b2?p9:b2))};
  assign y14 = (p0/a5);
  assign y15 = (!(a1|a4));
  assign y16 = (&($unsigned($signed((((p9!=p9)==(a0!=b1)))))));
  assign y17 = (-5'sd5);
endmodule
