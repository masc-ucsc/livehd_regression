module expression_00322(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~^(4'd9))==(~^(4'sd0)))?(((4'd4)*(4'sd3))<<((4'd7)<<<(3'd5))):(((2'd3)>>>(-2'sd1))*((2'd1)<=(3'd1))));
  localparam [4:0] p1 = ((3'd2)?(-2'sd0):(4'd6));
  localparam [5:0] p2 = ((4'sd6)!=(-4'sd5));
  localparam signed [3:0] p3 = (~^((~^(~(2'sd0)))<=(((5'd19)&&(3'd6))!=={4{(-2'sd1)}})));
  localparam signed [4:0] p4 = (-3'sd1);
  localparam signed [5:0] p5 = (((&(2'd3))>((3'd1)==(4'd11)))&(2'd2));
  localparam [3:0] p6 = (((-4'sd2)?(3'd7):(5'd17))?((3'd4)?(2'd2):(-4'sd0)):((3'd5)<=(5'd20)));
  localparam [4:0] p7 = {2{(4'd12)}};
  localparam [5:0] p8 = (({(5'd24),(-3'sd0)}?(!(5'd16)):(&(4'd3)))?(((-5'sd5)?(3'd6):(5'sd2))?((3'sd0)?(-4'sd1):(5'd17)):((3'd2)+(-4'sd6))):{(~&{{(4'd8),(2'd1),(-2'sd0)}})});
  localparam signed [3:0] p9 = (~^((|(((5'd12)?(5'd14):(4'd1))&((5'd8)?(-4'sd5):(2'sd1))))&&(((2'sd0)===(5'sd15))?((2'd1)>>>(4'd10)):(4'd2 * (5'd0)))));
  localparam signed [4:0] p10 = (({3{(-2'sd0)}}&&((2'd1)<(5'sd13)))==({4{(-4'sd4)}}^(-4'sd6)));
  localparam signed [5:0] p11 = ((!((3'd5)==(2'd3)))!=={(2'd0),(2'd0),(-5'sd15)});
  localparam [3:0] p12 = (((-5'sd15)<(3'd3))%(3'sd2));
  localparam [4:0] p13 = {2{{{{2{{(5'd24),(5'sd14),(4'sd0)}}}}}}};
  localparam [5:0] p14 = (((-3'sd1)?(2'sd1):(5'd28))?(!((5'd9)?(5'd17):(4'd6))):((-4'sd4)?(-3'sd1):(2'sd0)));
  localparam signed [3:0] p15 = {4{(!(|(|(5'd11))))}};
  localparam signed [4:0] p16 = {4{(!(4'd9))}};
  localparam signed [5:0] p17 = ({(-5'sd5),(3'sd0),(3'd1)}?((2'd0)?(-3'sd0):(5'd5)):{(3'd4),(2'd0)});

  assign y0 = (-2'sd0);
  assign y1 = (((((p7>=p14)||(p8))-((b4===a3)&(p9==p2))))>=$unsigned((($signed(p10)==(p5*p6))&((p15>p9)))));
  assign y2 = {($unsigned(((a3?a4:a3)))<=(5'd2 * $unsigned((b2))))};
  assign y3 = (({2{(|b2)}}>(b1?a1:p7))<<<({4{p13}}>>(~(p2?b0:p5))));
  assign y4 = (((~^(^(((a3-b1)^(~|a4))))))+$unsigned(((|(-a0))?(a0?b4:b3):(a3<<b1))));
  assign y5 = (b5|p9);
  assign y6 = (($signed((a2?a0:p13)))?(5'd2 * (p6|b2)):$unsigned(((b4===a4))));
  assign y7 = ($signed(({b4,a1,b3}!==(^b1)))?(!((p0)?(p16>=p13):(p13?p5:p12))):((p5?p14:p6)?(b2?p17:p1):(p0)));
  assign y8 = (~^($unsigned((p1))|((p5<=p0))));
  assign y9 = {($signed(b4)>>>{4{p2}}),{2{{3{b4}}}}};
  assign y10 = (((~^a4)?(a5/p16):(b2-b0))?(!((~&p1)?(^a4):(b5?p4:a1))):((^(2'd2))>>>(5'd5)));
  assign y11 = $unsigned((((~&$signed(p10)))?($unsigned((a1?a5:a2))):(!(!(+p6)))));
  assign y12 = {{(~|((&(&(~&$signed(a3))))=={(b3===b0),(a1&&p16),(^b0)}))}};
  assign y13 = ({{{3{b0}},(-p3)}}^{3{(b2?p0:a0)}});
  assign y14 = ((4'd12)>>>((p4>=p10)!=(b1?p3:a4)));
  assign y15 = {(((2'd1)>>>(5'd22))!=={(5'd7),(+a1),(a5-a0)})};
  assign y16 = (|((p6+p6)+(a2===b0)));
  assign y17 = $unsigned((($unsigned(p10)&&{1{b2}})!=$signed(($unsigned(a3)<(p8-b4)))));
endmodule
