module expression_00626(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({2{(-5'sd11)}}>(5'd11));
  localparam [4:0] p1 = (5'd2 * ((4'd10)!==(2'd1)));
  localparam [5:0] p2 = (|(2'd0));
  localparam signed [3:0] p3 = {3{(3'd3)}};
  localparam signed [4:0] p4 = (+(!(&(+(!((5'd5)<<<(3'd4)))))));
  localparam signed [5:0] p5 = (3'sd3);
  localparam [3:0] p6 = (((-((4'd7)>(2'd0)))|(^{((-5'sd8)>(3'd2))}))||((3'd3)!==(5'd25)));
  localparam [4:0] p7 = ((~^(~^((2'd0)<(2'd2))))<{{(-4'sd2),(5'sd1)},(~^(4'sd2))});
  localparam [5:0] p8 = (~&((-3'sd0)>>(4'd11)));
  localparam signed [3:0] p9 = (2'd1);
  localparam signed [4:0] p10 = ((4'sd3)^~(5'd4));
  localparam signed [5:0] p11 = (~&(+(|{(2'sd1),(4'sd5)})));
  localparam [3:0] p12 = (~&(~|{1{((((5'd6)-(4'd4))||((2'd0)&&(4'sd6)))>>>((+(4'd14))!=(!(4'sd3))))}}));
  localparam [4:0] p13 = {4{(3'd6)}};
  localparam [5:0] p14 = ((((5'sd8)&(-5'sd3))&((3'd7)<<(4'd3)))>={2{(5'd2 * (5'd1))}});
  localparam signed [3:0] p15 = ((((-2'sd1)?(-4'sd4):(-3'sd3))^~(2'd1))?((3'sd0)?(2'd3):(-4'sd2)):((2'd1)?(5'd31):(-2'sd1)));
  localparam signed [4:0] p16 = {3{(((-4'sd6)>(-2'sd0))=={(5'd10)})}};
  localparam signed [5:0] p17 = (((3'sd1)<<(2'd2))<=((-4'sd7)^(-4'sd1)));

  assign y0 = $unsigned({2{{2{(-p13)}}}});
  assign y1 = (4'd3);
  assign y2 = (($signed(p16)?(p9<p12):$signed(p7))?((b0)?{1{p14}}:(b2||a3)):({1{(b0>=a4)}}<=(p10^~b2)));
  assign y3 = (+(-$unsigned(p9)));
  assign y4 = {2{p2}};
  assign y5 = {({b3}?(6'd2 * b1):$signed(a0)),((a2>a2)<=(b3?a0:b1)),($unsigned((b5?a2:b2)))};
  assign y6 = (+(|((p17&&b0)<<(p12^~b2))));
  assign y7 = {((p17>=p10)<<(p3||p1)),({p3,p17,p12}-(~|p12)),((p8^~p16)|(a1^b4))};
  assign y8 = ((5'd2 * (p13&p6))<<((a0^p10)<(a2?p1:a0)));
  assign y9 = ((-5'sd14));
  assign y10 = (p11?p15:p14);
  assign y11 = (&(!{2{((|a4)?(a1?a1:a5):(~|a2))}}));
  assign y12 = (5'd14);
  assign y13 = (b5<b4);
  assign y14 = ({2{{1{b2}}}}>=((a4>>>b3)>{4{b5}}));
  assign y15 = {1{{2{(^{1{(p7&&p10)}})}}}};
  assign y16 = (2'sd1);
  assign y17 = {4{{3{a5}}}};
endmodule
