module expression_00413(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-3'sd2)||(4'd5));
  localparam [4:0] p1 = ((5'd2)<<(2'd3));
  localparam [5:0] p2 = ((^(!{(5'sd5),(-2'sd1),(5'd12)}))?(!(~^((3'sd0)<(-4'sd4)))):(~^{((-4'sd2)?(5'd18):(4'd10))}));
  localparam signed [3:0] p3 = (3'd4);
  localparam signed [4:0] p4 = ({1{(|((-2'sd0)?(3'sd1):(-4'sd2)))}}?((-3'sd2)?((2'd1)?(5'd17):(4'd5)):((-5'sd14)?(5'd16):(4'd14))):(!((-4'sd1)?(3'd1):(3'd3))));
  localparam signed [5:0] p5 = {(~(+(-{(5'd3),(2'd0)})))};
  localparam [3:0] p6 = ({3{{1{(-2'sd1)}}}}!={1{{2{{4{(5'd2)}}}}}});
  localparam [4:0] p7 = {3{(~^((~(5'd26))>>>(3'd4)))}};
  localparam [5:0] p8 = {1{({4{(3'sd1)}}?(4'sd3):(((5'd9)?(5'd24):(3'd5))?{3{(2'd2)}}:(2'd3)))}};
  localparam signed [3:0] p9 = ((5'd16)?(-2'sd0):(3'd5));
  localparam signed [4:0] p10 = (~|((^{((2'd2)>=(5'sd15)),{(~&(3'd4))}})!==(|{3{{2{(5'd5)}}}})));
  localparam signed [5:0] p11 = ((((-3'sd0)>>(4'd9))===((-2'sd1)+(-2'sd1)))?(((-4'sd3)^(-5'sd4))%(-2'sd0)):(((5'd14)&&(2'sd1))/(3'sd2)));
  localparam [3:0] p12 = {((4'd6)|(-2'sd0)),((3'd2)-(2'sd1))};
  localparam [4:0] p13 = (2'd0);
  localparam [5:0] p14 = (({(4'd3)}>={4{(3'sd2)}})?(+(!(-(~&(4'sd7))))):{{4{(3'd6)}}});
  localparam signed [3:0] p15 = (~&(!{{3{(+{(4'd7)})}}}));
  localparam signed [4:0] p16 = (((2'd1)>>(4'sd6))?((5'sd9)<<(2'd0)):((4'd12)==(2'd0)));
  localparam signed [5:0] p17 = ((((4'sd2)===(3'sd0))^((-2'sd1)!=(-5'sd9)))<<<(((-2'sd0)===(3'd2))&&{2{(4'sd6)}}));

  assign y0 = (!{4{(a5>>>b1)}});
  assign y1 = (|(({(~&(5'sd15))}<(3'd6))>({p12,b0,a3}<<<((&p14)!=(~b1)))));
  assign y2 = (((({b4}&&(b0===a4))^({4{p11}}<=(p16+a0)))>$unsigned({4{(p7&b4)}})));
  assign y3 = {4{({4{p3}}>{2{p16}})}};
  assign y4 = ((3'sd2)?(4'sd7):((a0&a2)<=(!(5'd15))));
  assign y5 = {4{{2{b1}}}};
  assign y6 = ((-$signed(($signed((p7?a4:a4))&((b5?b0:a5)))))>>(&(&((+{3{(p6?p8:a1)}})))));
  assign y7 = ((-(~|(5'd13)))!==(!({3{a3}}^~(4'd13))));
  assign y8 = ((-3'sd3)<=$signed(p2));
  assign y9 = (~&((-(p10?p17:p17))==(!(p4?p14:b3))));
  assign y10 = {((({p12,a0,p15}<(p4))!=((p15)+(p6?b5:p0)))&&{(!{p14,p10,a0}),$signed((b5|p17)),(p15>>>p11)})};
  assign y11 = {1{$signed((~^(($signed({2{p11}})<<<(p10^~p2))&(~|(-{3{{3{p15}}}})))))}};
  assign y12 = (((p1?p7:p7)>=($unsigned(p12)!=(p11>>>p14))));
  assign y13 = ((^(((+b3)>>(a1<<<b3))===(4'd11)))!==(6'd2 * (5'd2 * a1)));
  assign y14 = ({2{((p14<=p16))}}+((p6?p16:p6)?(p2>p2):(a4||p5)));
  assign y15 = (((b2?a3:a4)?(~^a3):(-a3))>((b2&&b1)>=(+b2)));
  assign y16 = (~^{1{((~(-{2{(-4'sd0)}}))^{3{(p3?p13:p13)}})}});
  assign y17 = (((b3?p4:p14)?{p13,p17,p17}:(p7?p16:p10))?({4{p3}}?(p6?p2:p3):(p8?p5:p15)):{{3{{3{p10}}}}});
endmodule
