module expression_00723(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((&(|{4{(4'sd4)}}))?{1{(2'sd1)}}:(-4'sd3));
  localparam [4:0] p1 = ((|(2'sd1))<<<((3'sd1)%(5'd5)));
  localparam [5:0] p2 = (-3'sd0);
  localparam signed [3:0] p3 = ((((-3'sd1)<=(2'sd0))!==((3'd5)<<<(4'sd6)))!=(((3'sd2)<=(-5'sd14))&((3'sd3)<(-3'sd3))));
  localparam signed [4:0] p4 = (3'sd3);
  localparam signed [5:0] p5 = ((((-3'sd0)^~(-3'sd2))>>((3'sd0)>>(5'd9)))|(((3'sd0)|(5'd15))-((4'sd6)>=(4'd6))));
  localparam [3:0] p6 = (((-2'sd0)?(4'sd4):(4'd15))?((5'd17)>(-4'sd3)):((4'sd1)>>(5'd20)));
  localparam [4:0] p7 = ({(5'sd10)}<((3'd0)-(5'd22)));
  localparam [5:0] p8 = (&(-(4'sd4)));
  localparam signed [3:0] p9 = (6'd2 * ((4'd5)<(3'd2)));
  localparam signed [4:0] p10 = (~({{(2'd1),(4'sd5)}}<<(^(~^(5'sd3)))));
  localparam signed [5:0] p11 = {{((2'd1)===(2'sd0)),{(3'd6),(5'd29),(3'd5)},{(-4'sd5),(3'd2)}},({(-5'sd0),(3'd6)}^~{(4'sd0),(3'd0)}),(4'd5)};
  localparam [3:0] p12 = {(2'd3),(3'sd2)};
  localparam [4:0] p13 = {(5'd12),(2'd1)};
  localparam [5:0] p14 = (^((5'd5)<=(3'sd0)));
  localparam signed [3:0] p15 = (+{(((4'sd0)&(4'sd1))^~(|((4'd14)?(4'd10):(-4'sd2))))});
  localparam signed [4:0] p16 = ((3'd3)>={1{(&{2{(2'd3)}})}});
  localparam signed [5:0] p17 = ((~^(5'd4))?((3'd6)!==(-5'sd8)):((5'sd6)?(5'd27):(4'd6)));

  assign y0 = (~&(5'd2 * {(+p1)}));
  assign y1 = ((((p5>>p9))<<<((p5>=p2)<<(p9>>b1))));
  assign y2 = (((2'd2)|(4'd6))^(5'd6));
  assign y3 = (4'd3);
  assign y4 = ($unsigned(($unsigned(p12)^(p3>=p1)))^{$unsigned(p16),(b3>=b1)});
  assign y5 = (((b4||b1)?(a1?b0:a5):(a0+b4))>={(~{(-{(a1>=a3),(b2?b3:p1),(b2+b4)})})});
  assign y6 = ((~|{2{({4{p16}}|(b4!=b4))}}));
  assign y7 = {{(p14||a3),(2'd2)},(3'd7),(-2'sd1)};
  assign y8 = (&(3'd4));
  assign y9 = (p16+p8);
  assign y10 = (p3?p17:p9);
  assign y11 = (((p7?p13:p10)+(~&(~&(p13?p8:p15))))>>((p7?p17:p3)?(~&(p7?p0:p3)):(p10?p17:p7)));
  assign y12 = {2{(b5>=p0)}};
  assign y13 = (!({4{(~|p1)}}?({2{p1}}>=(2'd1)):(3'd6)));
  assign y14 = (-{(b3+p11)});
  assign y15 = {2{{4{(a4?b4:p1)}}}};
  assign y16 = (|{(~&(a1!=b4)),((a5?b3:a2)-{a3,b0}),(-5'sd0)});
  assign y17 = {(a2!=b5),(^b1)};
endmodule
