module expression_00657(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&((4'd2)?((4'sd1)?(-4'sd4):(4'd9)):((4'd0)&&(5'sd8))));
  localparam [4:0] p1 = ({2{((5'd22)?(-4'sd5):(2'sd1))}}|(6'd2 * {1{{2{(3'd5)}}}}));
  localparam [5:0] p2 = ({(~(5'sd0)),(!(3'sd0)),(&(2'd3))}<(^{(4'd3),(2'd1),(2'd0)}));
  localparam signed [3:0] p3 = ((^{4{(5'sd6)}})?((-2'sd1)!==(3'sd2)):((5'd10)&&(3'd6)));
  localparam signed [4:0] p4 = (5'd2 * (5'd15));
  localparam signed [5:0] p5 = ({2{{(-3'sd1),(-2'sd0),(-3'sd0)}}}&{((2'd3)>>>(2'sd1)),((5'd22)^~(3'd5)),((4'd10)>>(2'd2))});
  localparam [3:0] p6 = (((5'sd14)?(4'sd4):(3'sd3))?((3'd0)?(3'd6):(4'd9)):((4'd4)?(-4'sd6):(2'sd0)));
  localparam [4:0] p7 = (~|(((5'sd14)>>(5'd24))>>((5'd12)<(2'sd1))));
  localparam [5:0] p8 = ((-(~^{((-4'sd7)?(3'd2):(3'd6))}))^(~|(((5'd24)<<<(-4'sd0))?(-(2'd1)):(!(-4'sd4)))));
  localparam signed [3:0] p9 = (+{((-2'sd0)?(3'd1):(-5'sd7)),(~|((5'd10)!==(2'd0))),((4'sd6)?(4'd15):(3'sd0))});
  localparam signed [4:0] p10 = (({2{(5'd3)}}!=((2'd0)===(2'd2)))<<{3{((5'd2)&(5'd10))}});
  localparam signed [5:0] p11 = ((4'd9)+((4'd7)?(3'd1):(5'sd0)));
  localparam [3:0] p12 = (~^{1{{3{((-5'sd5)^(2'd0))}}}});
  localparam [4:0] p13 = {3{(-4'sd1)}};
  localparam [5:0] p14 = (((-2'sd0)&&(2'sd1))?{3{(4'sd7)}}:((5'd31)>>(4'sd0)));
  localparam signed [3:0] p15 = ((-2'sd0)===(3'sd0));
  localparam signed [4:0] p16 = {1{(2'sd0)}};
  localparam signed [5:0] p17 = (((4'sd3)?(2'sd1):(-5'sd1))?((~^(2'sd1))>(-2'sd1)):(!{4{(5'd19)}}));

  assign y0 = (~^{2{p12}});
  assign y1 = (+{2{(+(~|{1{((&(b0!==a4))||(|(a4<a0)))}}))}});
  assign y2 = (~|{1{(^{1{{2{((p13||p8)^(^$unsigned(p11)))}}}})}});
  assign y3 = (^{(!(~^{p14,a2,a0})),(^(p8-a5)),(+{{p1,b0}})});
  assign y4 = (~^(+{{{p13}},(~{p10,p5}),{p6,p0}}));
  assign y5 = {3{((b5?p7:a4)>={3{p2}})}};
  assign y6 = {1{(~{1{(~&{2{{3{{2{p17}}}}}})}})}};
  assign y7 = {4{(a2?a1:b5)}};
  assign y8 = (^(b3!==a3));
  assign y9 = (~&{(+{((^{p14,b2,b5})?(b4?b0:b1):(a3?b1:b2))}),{((a1?a1:a5)>>(|(a2>>a2)))}});
  assign y10 = (((p10?p17:p14)|(b5!==a0))>>$signed((5'd2 * (p6<<p14))));
  assign y11 = $signed($signed((3'sd1)));
  assign y12 = (+(~|p5));
  assign y13 = {4{(!b5)}};
  assign y14 = ((^(~^{3{(a2&&b2)}}))!==(&{4{$unsigned(b4)}}));
  assign y15 = (~&(~^p3));
  assign y16 = (p1?p10:p17);
  assign y17 = $unsigned((&(4'd0)));
endmodule
