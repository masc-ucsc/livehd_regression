module expression_00539(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd7)<(5'd29));
  localparam [4:0] p1 = (((3'sd0)<=(3'd1))%(4'd5));
  localparam [5:0] p2 = {((2'd1)==(3'd2)),{((4'd11)==(-4'sd3))}};
  localparam signed [3:0] p3 = ({3{(5'd30)}}!==(&(3'd7)));
  localparam signed [4:0] p4 = {(|(&(5'sd13))),{(5'd3),(5'd29),(-2'sd1)}};
  localparam signed [5:0] p5 = ((4'd7)&&(((2'sd1)&(4'd1))^~(~|(2'd0))));
  localparam [3:0] p6 = {1{(6'd2 * (-((5'd6)+(3'd5))))}};
  localparam [4:0] p7 = ((-5'sd8)!==(5'd18));
  localparam [5:0] p8 = (+((&((-(5'd2))&&((5'sd6)^~(2'd3))))!=(((5'sd15)!==(5'd23))-((-5'sd0)%(3'sd1)))));
  localparam signed [3:0] p9 = (({2{(-4'sd7)}}<<((4'sd3)<(2'sd1)))>>(((5'd16)>=(-4'sd3))>(4'sd6)));
  localparam signed [4:0] p10 = (((3'd2)<(2'd3))?((4'd14)!==(-4'sd0)):{4{(5'sd14)}});
  localparam signed [5:0] p11 = (~((5'd28)>=(|(~(2'd1)))));
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = (!(((5'd26)<<<(3'd6))+{(4'd0),(-4'sd0)}));
  localparam [5:0] p14 = ((((2'd1)&&(2'sd1))||{2{(-2'sd1)}})<(~&((4'd14)>=(3'd6))));
  localparam signed [3:0] p15 = {(-2'sd0)};
  localparam signed [4:0] p16 = ((!(+(3'd4)))/(2'd2));
  localparam signed [5:0] p17 = ((!(5'd28))?((-4'sd1)?(2'sd1):(3'sd2)):(^(3'd4)));

  assign y0 = (~(((p16>>>b4)<(a3-p3))<(~^(~&(a4<<<p6)))));
  assign y1 = {($signed(((b3?p3:p6)?(b1?b0:b4):$unsigned(p7)))?$unsigned(((a5!==b2)&&(b3-b3))):((p2<=b2)?(p3):{2{p7}}))};
  assign y2 = ((~(~|a3))<<<(p6||p17));
  assign y3 = ((!((p17+b3)&{p12,p7}))<((b3<=a0)>{p14,a2,a5}));
  assign y4 = (3'd1);
  assign y5 = (~^(((!$unsigned(p6))>>(p7<<<a5))>>((~|$signed(b0))<=(p12>>p11))));
  assign y6 = ((4'd15)<<<(~(|p0)));
  assign y7 = (~(^((~^p0)>(+a3))));
  assign y8 = (~|((&{(4'd10),(p16<<<p2),(b1===a2)})>>((5'd21)-((-5'sd11)^~(!p10)))));
  assign y9 = {(-3'sd3),((a4||b1)&(2'd0)),(^((b5<<a5)?(-3'sd3):{a2}))};
  assign y10 = (((~(^a0))>>>(|(^b4)))?((!p5)?(~|b4):(^a0)):(~|{(~&b0),(b4||b2)}));
  assign y11 = ({4{p12}}>>>(!(^b4)));
  assign y12 = (~^(+(|p16)));
  assign y13 = (~|(~^{4{(3'd5)}}));
  assign y14 = ((p13?p1:p13)+(p8>>>p17));
  assign y15 = ((2'd2)<<<((^(-3'sd2))!==(|(-a0))));
  assign y16 = {2{$signed({1{{3{{4{a0}}}}}})}};
  assign y17 = $unsigned((5'sd13));
endmodule
