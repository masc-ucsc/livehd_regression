module expression_00222(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{((-2'sd1)^(-2'sd1))}}+{4{{(4'sd1)}}});
  localparam [4:0] p1 = {((5'd27)?(4'd12):(-5'sd7)),(|(2'sd0))};
  localparam [5:0] p2 = {2{{4{(3'd0)}}}};
  localparam signed [3:0] p3 = (~(((~&(5'd3))?(~^(3'sd3)):((4'sd0)<<<(-4'sd6)))==(^(~&(((2'd1)<<(2'd3))>>{2{(-4'sd7)}})))));
  localparam signed [4:0] p4 = {1{(-5'sd4)}};
  localparam signed [5:0] p5 = {1{{1{({4{(3'd6)}}+({3{(3'd4)}}<<((-2'sd0)<(3'sd2))))}}}};
  localparam [3:0] p6 = (((3'd7)>>(3'sd0))<<((-2'sd0)%(-3'sd2)));
  localparam [4:0] p7 = ((!(4'd14))>>>((5'd8)==(-5'sd5)));
  localparam [5:0] p8 = (!(3'd0));
  localparam signed [3:0] p9 = (((5'sd10)>>>(4'sd5))>>>((-2'sd1)?(2'd1):(5'd0)));
  localparam signed [4:0] p10 = (((3'd0)!=(-3'sd3))<((-3'sd1)!=(5'd3)));
  localparam signed [5:0] p11 = (((-2'sd0)|(3'd6))^(-(-2'sd1)));
  localparam [3:0] p12 = (3'd2);
  localparam [4:0] p13 = (5'd0);
  localparam [5:0] p14 = {4{(5'd5)}};
  localparam signed [3:0] p15 = (+(!(((2'd0)?(4'sd2):(4'd13))?((2'd0)<<<(-3'sd3)):((2'd0)?(2'd2):(-5'sd15)))));
  localparam signed [4:0] p16 = (2'sd1);
  localparam signed [5:0] p17 = {3{{(-4'sd7),(2'd2)}}};

  assign y0 = (({p2,p1,p17}&&(!{a3,p6}))^(5'd2 * (~&$unsigned(a3))));
  assign y1 = (((|(!a3))<(~(b5>=a0)))!=(~({a1,a1}!==(b1==a3))));
  assign y2 = ((p14+a1)?(~{b1,a1,b5}):$signed((p8?b5:b0)));
  assign y3 = (!(~{2{a5}}));
  assign y4 = (5'd20);
  assign y5 = (a1^~a5);
  assign y6 = {2{((&($unsigned($signed(b1)))))}};
  assign y7 = (+((&(2'd1))?{p12,a1,b4}:(5'sd15)));
  assign y8 = (~^(^(+{p1})));
  assign y9 = (((^a2)*(|a1)));
  assign y10 = ((4'd13)||{4{{2{p13}}}});
  assign y11 = {4{(~^p15)}};
  assign y12 = ((5'd9)<{{p10,p10,p12},(p16)});
  assign y13 = (-4'sd5);
  assign y14 = (-5'sd0);
  assign y15 = ({1{(5'sd2)}}?({1{p3}}?{1{a3}}:(b3?p17:p9)):{2{(3'd7)}});
  assign y16 = ({2{(~|({1{p9}}!=(p1<p15)))}}^~(|{3{(~(p3^p17))}}));
  assign y17 = ((a3-b5)&&(a3==a4));
endmodule
