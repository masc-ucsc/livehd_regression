module expression_00129(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'd0)?(2'sd1):(5'sd1))?{3{(5'd7)}}:(|(2'd0)))?((&(3'sd1))?{3{(5'd29)}}:{2{(5'sd10)}}):(((4'd15)?(3'd5):(5'd7))?((3'd1)?(3'sd0):(5'd11)):(+(5'sd11))));
  localparam [4:0] p1 = (-(&(4'd9)));
  localparam [5:0] p2 = {(((-2'sd1)?(2'd2):(5'd27))?(6'd2 * (2'd0)):((-2'sd0)?(2'd2):(-4'sd5)))};
  localparam signed [3:0] p3 = (-(~{3{(+(|(-3'sd2)))}}));
  localparam signed [4:0] p4 = (~&(((-2'sd0)&(2'sd1))<<<((3'd0)?(-5'sd0):(3'sd2))));
  localparam signed [5:0] p5 = ((((-5'sd9)!==(5'd1))?(-3'sd0):{3{(3'd2)}})?((~^(4'd6))?{4{(2'sd1)}}:(2'sd0)):(3'd4));
  localparam [3:0] p6 = (2'd0);
  localparam [4:0] p7 = (~|(!((!{1{(+(~|{1{(-4'sd6)}}))}})^~({2{(4'd3)}}<<{3{(3'd0)}}))));
  localparam [5:0] p8 = ((+(4'd1))>=(~|(-4'sd6)));
  localparam signed [3:0] p9 = (3'd7);
  localparam signed [4:0] p10 = (3'sd2);
  localparam signed [5:0] p11 = (&(((2'd0)||(3'd0))>>>(((5'd28)<<(3'sd1))!==(~&{(-2'sd1),(4'd2)}))));
  localparam [3:0] p12 = (+(((4'd13)?(-3'sd0):(5'sd1))!={4{(-5'sd6)}}));
  localparam [4:0] p13 = ((((4'd9)?(5'd7):(3'd2))?((2'd1)>(3'd2)):{(5'sd9),(5'sd2)})>>>(((-4'sd1)&(4'd0))<={3{(-3'sd3)}}));
  localparam [5:0] p14 = (((2'd1)?(4'd4):(3'd6))^(((3'd0)?(5'd31):(3'd6))>((-3'sd3)?(5'd19):(3'sd0))));
  localparam signed [3:0] p15 = (~((4'd6)<<<(2'sd0)));
  localparam signed [4:0] p16 = (((2'd3)!=(4'd0))==((2'sd1)|(2'd2)));
  localparam signed [5:0] p17 = (&(~&(~|(-((!(&(~(-4'sd0))))!=((~&(4'sd5))>>(3'd4)))))));

  assign y0 = $signed($unsigned((p13?p17:p4)));
  assign y1 = (~|(~((~|(~&(-$unsigned((~(~|$signed((&((&p0)||(+a1)))))))))))));
  assign y2 = ($unsigned(p0)?(b2<=p7):(p6?b5:b1));
  assign y3 = (!(~&(p14<<p12)));
  assign y4 = {2{{1{(3'd4)}}}};
  assign y5 = ((4'sd6)?(-3'sd1):(5'd2));
  assign y6 = $unsigned(((2'd3)|((p0?p0:b0)|(~^(^p3)))));
  assign y7 = $signed({{3{$signed(b3)}},{{3{a0}}},{2{(2'd1)}}});
  assign y8 = ((+b3)<(~|p10));
  assign y9 = ((((-a5)||(~^b1))<<((p0?p5:a4)-(&p12)))<<(+($unsigned(((b3)))>>>(^(b0-b2)))));
  assign y10 = (({1{{(p9>=p15)}}}^{3{{1{a1}}}})-(((a0>>>p13)||{p17,p8,p10})||({1{p17}}^~{p17,b4})));
  assign y11 = (~&(~{{(~^p0),{p10}},({p2}!=(+a4))}));
  assign y12 = ((((^a5)==(a2>=b5))&$signed((a3^~b3)))!==(^$signed($unsigned((^(b2?a0:a3))))));
  assign y13 = (4'd9);
  assign y14 = (-2'sd0);
  assign y15 = ({(a3?p15:p13),{a5,p1}}&&{(|p3),$signed(p3),{1{a5}}});
  assign y16 = (!{{(&({(-{a0,p10,a0})}<=(3'd4)))}});
  assign y17 = (5'd2 * b2);
endmodule
