module expression_00120(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd11);
  localparam [4:0] p1 = {{{{(-2'sd1),(4'd1)},{(4'd15)},{(3'sd3),(5'd17)}},{{{(3'sd1)},{(5'd27),(3'd1),(4'sd7)}}},{{(2'sd0),(3'd2),(4'sd4)},{(3'sd1)},{(2'd0),(-5'sd14),(5'd8)}}}};
  localparam [5:0] p2 = (5'd11);
  localparam signed [3:0] p3 = ((5'd23)!=(5'sd1));
  localparam signed [4:0] p4 = ((((4'd2)&&(-5'sd7))?{2{(3'd3)}}:((-3'sd3)+(2'sd0)))===(((5'd22)?(-2'sd1):(-5'sd2))>>>((3'd7)>>(5'd23))));
  localparam signed [5:0] p5 = {4{((5'd24)?(-2'sd0):(5'sd14))}};
  localparam [3:0] p6 = (~&{4{{1{((-2'sd0)?(4'd4):(2'd3))}}}});
  localparam [4:0] p7 = {4{(5'sd15)}};
  localparam [5:0] p8 = (~|{4{(-(5'd30))}});
  localparam signed [3:0] p9 = (3'd1);
  localparam signed [4:0] p10 = ({3{{2{(3'sd3)}}}}?{2{((4'd8)>(-2'sd1))}}:({3{(4'd4)}}=={2{(5'd21)}}));
  localparam signed [5:0] p11 = ((((5'd12)>(3'd2))>>((2'd2)<(5'sd2)))>>>(4'd2 * (5'd2 * (4'd10))));
  localparam [3:0] p12 = (~^(+{2{(-2'sd0)}}));
  localparam [4:0] p13 = {1{{1{{3{{1{{3{(-4'sd2)}}}}}}}}}};
  localparam [5:0] p14 = ({3{((2'd1)<(-2'sd1))}}-(-((~^((2'sd0)<<<(4'd0)))===(&(+(5'd6))))));
  localparam signed [3:0] p15 = {{{(-2'sd1),(3'd5),(2'd0)},{(5'sd6)},(&(-2'sd0))}};
  localparam signed [4:0] p16 = ((((2'd0)?(5'sd6):(-2'sd1))/(-3'sd2))&&(((2'd1)/(5'd13))?((5'd19)<=(2'd3)):((2'd3)%(5'sd12))));
  localparam signed [5:0] p17 = ((-4'sd2)|(4'd3));

  assign y0 = ({2{p3}}&&(p15^b5));
  assign y1 = (b1+a3);
  assign y2 = (-4'sd1);
  assign y3 = (b1?a3:a5);
  assign y4 = $signed((-((|{4{{1{p11}}}})&&(+(!($unsigned(p3)?(~^p5):{4{p13}}))))));
  assign y5 = (((&b1)?$signed(a5):(-b2))?{(a2<=b2),(a0<b5)}:((!$unsigned(a3))!=={b2,b4}));
  assign y6 = ((a5|p2)!={2{a4}});
  assign y7 = ({(p1?p16:p6),(p9?p6:p12),(p15?p11:b3)}?((a2?p6:p11)+(a0?a2:p4)):{(a1===b0),(!p4),{p16,p7}});
  assign y8 = {a2,p10,b3};
  assign y9 = (($unsigned(p6)?{a3}:(p1?p9:p17))?((~|p9)&&(p0)):({p12}?(p12-p3):{p0,p2,p1}));
  assign y10 = ({1{{4{(a2>b2)}}}}>=(^(~&(^((6'd2 * b1)<<<(-a0))))));
  assign y11 = ((^(p15?p9:p4))>>>(~|({p14,p10,p12})));
  assign y12 = (4'sd5);
  assign y13 = (2'sd0);
  assign y14 = ((3'd7)||(((a3?a1:a5)?(4'd10):(-3'sd1))<(-5'sd12)));
  assign y15 = (2'sd0);
  assign y16 = (($signed(((~^{3{(b3?a3:a1)}})))));
  assign y17 = (p15<=p6);
endmodule
