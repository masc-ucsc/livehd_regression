module expression_00299(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(&((&(~|(&((5'd27)==(5'd17)))))>=((~&(-3'sd0))<<<((4'd13)<<(-3'sd3))))));
  localparam [4:0] p1 = ((~(-(!(~(-((2'sd0)&(5'sd0)))))))>((+((5'd25)<<(4'd4)))<<<(((2'd0)/(-2'sd1))+(~^(3'sd1)))));
  localparam [5:0] p2 = {(((-3'sd1)?(2'd1):(3'd7))?(-2'sd0):{(5'sd2),(2'd2)})};
  localparam signed [3:0] p3 = (~(+(((2'd1)?((3'sd3)&(-2'sd1)):(|(-2'sd1)))>>(((4'd10)>=(5'sd7))-(&(4'sd7))))));
  localparam signed [4:0] p4 = ((((5'sd8)>=(4'd9))>>((3'sd0)+(-5'sd5)))>(|(!((-5'sd7)>>(5'd20)))));
  localparam signed [5:0] p5 = (2'd2);
  localparam [3:0] p6 = (((3'd3)?(-5'sd9):(-4'sd1))?{2{(3'd4)}}:((-2'sd1)>>>(-2'sd0)));
  localparam [4:0] p7 = ({4{(2'd0)}}<((4'd5)>>>(-3'sd0)));
  localparam [5:0] p8 = ((&(|((5'sd10)||(2'd3))))>=((5'd22)?(2'sd0):(4'sd0)));
  localparam signed [3:0] p9 = (+(+(^(~&(~{4{(|(!(3'd2)))}})))));
  localparam signed [4:0] p10 = ({1{((^(4'sd7))===((4'd9)&(5'd6)))}}&(+{3{(-3'sd2)}}));
  localparam signed [5:0] p11 = ((((-4'sd7)?(2'sd1):(2'd0))?{(-3'sd1)}:(-(-3'sd1)))?({(2'd0)}+(~&(-2'sd1))):(((4'sd5)<<<(5'd6))?((4'd3)?(-3'sd2):(4'd12)):(|(3'd2))));
  localparam [3:0] p12 = (|(|(+(3'd1))));
  localparam [4:0] p13 = ((((5'd1)?(5'sd1):(3'd5))||(~|((-3'sd1)!=(2'd3))))|((|((5'sd6)?(3'sd0):(2'sd0)))>((4'd10)?(2'd2):(2'd0))));
  localparam [5:0] p14 = (2'd2);
  localparam signed [3:0] p15 = (&(-5'sd14));
  localparam signed [4:0] p16 = {{(3'd4),(5'd12),(3'd4)},((4'd13)?(3'd0):(2'd2)),(3'sd0)};
  localparam signed [5:0] p17 = (~|((((3'sd3)==(-3'sd2))&&((5'd16)>=(3'sd1)))>>(((5'd11)|(-2'sd0))?((3'd6)?(2'd2):(5'd29)):((3'd7)==(5'd0)))));

  assign y0 = (^(!{2{(^(&(~^((~&p8)))))}}));
  assign y1 = $signed(p13);
  assign y2 = (+((p6||a3)?(p8?p17:a2):(~&(p16+p9))));
  assign y3 = {$unsigned((~{3{{1{p10}}}})),{{b3,p17},$unsigned(p16),{a3,p1,p11}},{{p15,p5,p5},$signed({p8})}};
  assign y4 = (a2?b2:b3);
  assign y5 = ((~&$signed({4{p14}}))=={3{$unsigned(p14)}});
  assign y6 = ((&(^((p3<=p7)&(-b3))))+((^{b4,a2})!=={{b2}}));
  assign y7 = (~&(!(!(2'sd0))));
  assign y8 = (-2'sd1);
  assign y9 = (^(~&(~&((~&((^p7)?(~&p2):(~&p1)))?((+(~&p13))<=(p14&a3)):{(+(~^a5)),(~&{p1,p1,p12})}))));
  assign y10 = {3{{4{{2{b2}}}}}};
  assign y11 = (p12+p0);
  assign y12 = (6'd2 * (p1?b0:b1));
  assign y13 = (~((|b5)&&{1{p11}}));
  assign y14 = $unsigned((3'd5));
  assign y15 = {2{(4'd0)}};
  assign y16 = (((~p0)?(p2|b1):(p16?p4:a4))<<((a4&p12)?(p16==p3):(b0<p9)));
  assign y17 = $unsigned({3{{2{(p17&&p11)}}}});
endmodule
