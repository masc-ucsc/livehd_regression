module expression_00489(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-3'sd2)?(5'd3):(2'sd0))>>((3'sd0)<<<(-5'sd4)));
  localparam [4:0] p1 = {2{({4{(5'sd13)}}^((-4'sd2)===(-4'sd4)))}};
  localparam [5:0] p2 = (!(4'd0));
  localparam signed [3:0] p3 = (((4'd14)?(5'sd5):(5'd3))?((3'd0)?(-3'sd3):(-3'sd2)):((5'sd12)?(-4'sd2):(4'sd3)));
  localparam signed [4:0] p4 = (~|(-4'sd6));
  localparam signed [5:0] p5 = ((-5'sd7)^(5'sd5));
  localparam [3:0] p6 = ((3'sd0)>((5'sd6)?(3'd1):(4'sd0)));
  localparam [4:0] p7 = {2{(6'd2 * (+(5'd17)))}};
  localparam [5:0] p8 = ((((5'sd8)^~(-2'sd0))?((2'd0)?(4'sd2):(3'd1)):{3{(-4'sd2)}})||({(2'd0),(-2'sd1)}<<{3{(5'd28)}}));
  localparam signed [3:0] p9 = ((((-5'sd7)>(5'd13))-((-4'sd5)<=(-5'sd9)))<(((-2'sd1)==(2'd0))^((-3'sd3)===(5'd2))));
  localparam signed [4:0] p10 = (^(((3'd0)==(-4'sd1))?((2'd0)!=(-5'sd9)):{(4'd15)}));
  localparam signed [5:0] p11 = (3'd6);
  localparam [3:0] p12 = (~^{(5'd17)});
  localparam [4:0] p13 = ({(-4'sd3)}=={1{(2'd0)}});
  localparam [5:0] p14 = (-4'sd2);
  localparam signed [3:0] p15 = (^((((2'sd0)?(5'd15):(-4'sd2))<<<((3'sd3)&(3'sd2)))?(~&((4'sd5)?(3'sd0):(2'd0))):((5'd14)?(3'sd3):(5'd4))));
  localparam signed [4:0] p16 = (&{3{{2{(3'd0)}}}});
  localparam signed [5:0] p17 = (-{3{(&{2{(5'sd5)}})}});

  assign y0 = (a4&&p5);
  assign y1 = (!(5'd2 * {1{(~&b0)}}));
  assign y2 = {2{p14}};
  assign y3 = (-(~|((-b4)<<<(~^a5))));
  assign y4 = (~|(~(^(&(~^(!(~(~&(~|(~&(~|(^b3))))))))))));
  assign y5 = (a4?a5:b3);
  assign y6 = ((p16|p0)<<{4{p6}});
  assign y7 = (a5|p13);
  assign y8 = (!(&{4{(4'd15)}}));
  assign y9 = ({2{a4}}<<<(a5!==a2));
  assign y10 = (((a4+b4)<<<(a4&a2))||((p6%a0)&(b5>b0)));
  assign y11 = (5'd21);
  assign y12 = $unsigned((5'd24));
  assign y13 = (((a4?p15:p14)?$signed($unsigned($signed(p6))):$unsigned((p7?p0:p12))));
  assign y14 = ((a5<=a0)!==(b0>>b4));
  assign y15 = ($unsigned(($unsigned($unsigned(a1))>>{a0,p17,p4}))!={(p11&b2),(a4!=p17),$unsigned(p0)});
  assign y16 = ((&{1{((~^(b1^~b1))!==(a1<<<b1))}})^(&(+(^(-(|(a2?b3:p2)))))));
  assign y17 = {((p9&&a1)&&(|$unsigned(p8))),{{2{p0}},$unsigned(a1),(~&p3)},(((-(b5===a2))<<<((p3!=a2))))};
endmodule
