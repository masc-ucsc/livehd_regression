module expression_00757(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd3);
  localparam [4:0] p1 = (+((-5'sd9)&&(!(((4'd3)>=(4'd5))+((2'd0)+(4'd13))))));
  localparam [5:0] p2 = {(3'd1),(4'sd1),(4'd15)};
  localparam signed [3:0] p3 = ((((2'd3)||(2'sd0))!==((4'd2)+(2'd1)))||(((3'sd1)<=(5'sd0))%(-5'sd0)));
  localparam signed [4:0] p4 = ((-4'sd0)^~(-3'sd0));
  localparam signed [5:0] p5 = (((3'd6)&&(-2'sd0))*(4'sd7));
  localparam [3:0] p6 = (^{((-3'sd1)<<<(4'd15))});
  localparam [4:0] p7 = ((5'd5)===(4'd15));
  localparam [5:0] p8 = (5'sd0);
  localparam signed [3:0] p9 = {1{(((2'd2)^~(2'sd0))?((3'sd3)?(4'd6):(5'd24)):((2'sd1)>=(4'sd2)))}};
  localparam signed [4:0] p10 = (3'd7);
  localparam signed [5:0] p11 = (((-3'sd1)?(3'd0):(5'd23))?{((3'd0)?(3'd6):(4'd8))}:((-4'sd7)?(-2'sd1):(5'd13)));
  localparam [3:0] p12 = ({{(2'sd0),(5'd2 * (3'd4)),(4'sd4)}}+{(|((-4'sd4)>>>{(4'd0),(4'd11),(4'd3)}))});
  localparam [4:0] p13 = (~|(~^{4{(4'sd3)}}));
  localparam [5:0] p14 = ((3'sd0)^((2'd2)^(4'd7)));
  localparam signed [3:0] p15 = (((-2'sd1)>>(|(3'd5)))<={2{(!(4'sd1))}});
  localparam signed [4:0] p16 = (3'd4);
  localparam signed [5:0] p17 = (^(&((-(3'sd1))?((5'd5)?(-3'sd3):(-4'sd2)):((-5'sd6)?(2'd2):(5'sd10)))));

  assign y0 = ((4'd2 * $unsigned((b0<=p7)))!=$signed(({a3,b0})));
  assign y1 = ({2{(p6?p8:b4)}});
  assign y2 = {(~&(5'sd10)),((b5?b3:b3)<=(a3?a5:b3)),((b1||a3)>>>(a2?b5:a5))};
  assign y3 = (!({3{(a4^~a4)}}?((&((b4)!=={b1}))):((-2'sd0)?(+a1):(b5?a4:b0))));
  assign y4 = {({(b4<=b4),(b2==a0),{1{a3}}}>={3{{2{a1}}}})};
  assign y5 = (^(((3'd7)?(+p0):(~&p10))&&(5'sd6)));
  assign y6 = (!{(+(!{p13,p15,p1})),(5'd18),(5'd31)});
  assign y7 = {p4,a1};
  assign y8 = $unsigned($unsigned($signed((5'd2 * $unsigned((5'd2 * p2))))));
  assign y9 = ({{p11},(-2'sd0),(p16^~p6)}-{2{(4'sd6)}});
  assign y10 = (+(&(&(^p13))));
  assign y11 = (+(~&((p5^p11)||$unsigned((p4==p14)))));
  assign y12 = (~^(p17||p1));
  assign y13 = (&(+(p0>=p13)));
  assign y14 = {4{(~&(~^(&p15)))}};
  assign y15 = (-$signed((~|(~^($unsigned((((~^b4)|$signed(p8))))<=(~&(~^(-2'sd1))))))));
  assign y16 = (5'd14);
  assign y17 = ((!(~^(|(4'd13))))&&((2'd1)>>(&(-5'sd13))));
endmodule
