module expression_00410(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd13);
  localparam [4:0] p1 = {1{(4'sd6)}};
  localparam [5:0] p2 = ((~&{(3'd1),(5'd29)})^{(-5'sd5),(-5'sd7)});
  localparam signed [3:0] p3 = ((((4'd1)===(2'd0))/(-4'sd6))-((4'sd4)?(4'd12):(-3'sd3)));
  localparam signed [4:0] p4 = (!(&{((5'd3)||(2'sd1)),{(5'd4),(2'sd0),(-2'sd0)},(&(2'd3))}));
  localparam signed [5:0] p5 = (~&(-2'sd0));
  localparam [3:0] p6 = (&((~(~|(!((3'd3)>(-5'sd3)))))&(((2'd3)^(3'sd2))>>(~^(~|(4'd13))))));
  localparam [4:0] p7 = ((~(|(!(4'sd2))))<<<((~|(4'sd5))<=(|(2'd1))));
  localparam [5:0] p8 = {(((3'd0)?(3'd6):(5'sd6))&(2'd3)),({(2'd1)}?((-3'sd2)?(5'sd5):(2'd0)):(3'd4))};
  localparam signed [3:0] p9 = {3{{1{((2'd3)<=(-5'sd11))}}}};
  localparam signed [4:0] p10 = (-((4'd10)?(-3'sd0):(2'd3)));
  localparam signed [5:0] p11 = (~(3'd2));
  localparam [3:0] p12 = {({{(2'd2),(-2'sd1),(2'd3)},(5'd27)}<=(((5'd29)<<(4'd14))!=((-2'sd1)&&(2'd0))))};
  localparam [4:0] p13 = (((5'd6)|(4'sd3))<=((3'd4)||(3'd2)));
  localparam [5:0] p14 = (~((4'd7)/(4'd13)));
  localparam signed [3:0] p15 = (|((~{(-3'sd2)})!=={{(-4'sd3),(3'd1)}}));
  localparam signed [4:0] p16 = (|(3'd7));
  localparam signed [5:0] p17 = (5'd23);

  assign y0 = (5'd2 * (b0>>p8));
  assign y1 = (~&(^(((b2==a5)>>(3'sd0))^$unsigned((-4'sd1)))));
  assign y2 = (p11<<<p1);
  assign y3 = ({4{b2}}?(b1?p8:p16):(&$unsigned(a0)));
  assign y4 = ((~^(~^(a2<b1)))!==$signed((-(~(a4*a2)))));
  assign y5 = $signed(((b2>=a3)?(p13):(|p0)));
  assign y6 = ({1{(p9<<p10)}}<<{4{p2}});
  assign y7 = ((~&(&b4))>=(b5>=p5));
  assign y8 = ({4{a1}}<<(~^((~|p14)>>(!b0))));
  assign y9 = {(p5>>b4),(p9?a4:p15),(a0?p11:a5)};
  assign y10 = (!(|(~&((p16&&p3)&{4{p5}}))));
  assign y11 = (^((p3?a5:a3)?(b3||p8):(~(b2?b1:p10))));
  assign y12 = (+(&((&(~&((^b2)>>(a5<b5))))!=$unsigned($signed((~(^(a2<b3))))))));
  assign y13 = {3{(3'sd0)}};
  assign y14 = ({3{(b1==b0)}}|(5'sd13));
  assign y15 = (($signed(p0)?(b5!==a3):(-p7))?$signed({{p11},(p11<p5)}):($signed(b3)?(p10-p7):$signed(b1)));
  assign y16 = ($signed((~^(-2'sd0)))?(2'd1):((~&a0)?(|b3):(b0)));
  assign y17 = (5'd1);
endmodule
