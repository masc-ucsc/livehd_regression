module expression_00067(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(~^(((3'd4)?(-3'sd1):(3'sd2))?{(!(3'sd0))}:(!{(4'd7)}))));
  localparam [4:0] p1 = (2'sd0);
  localparam [5:0] p2 = ((2'sd0)^(5'd11));
  localparam signed [3:0] p3 = (-3'sd0);
  localparam signed [4:0] p4 = (5'd2 * {(2'd3),(2'd1),(2'd1)});
  localparam signed [5:0] p5 = (((-3'sd1)?(3'd3):(3'd1))-((-2'sd1)?(-2'sd1):(4'd3)));
  localparam [3:0] p6 = (^((~|(3'sd2))&(-2'sd1)));
  localparam [4:0] p7 = {(~|((5'd7)?(5'sd9):(4'sd2))),((3'd7)?(-2'sd0):(-3'sd3))};
  localparam [5:0] p8 = {({(5'd6),(4'sd6),(2'd2)}>={(5'd28),(2'sd1),(4'd6)})};
  localparam signed [3:0] p9 = (|((((-2'sd1)-(-3'sd2))!=((2'd3)|(5'd2)))!=((^(2'd1))*((5'd9)<<<(2'd3)))));
  localparam signed [4:0] p10 = (2'd1);
  localparam signed [5:0] p11 = (((-2'sd0)^~((3'd0)==(2'd0)))|({4{(5'd13)}}?(2'd2):((-2'sd0)?(5'sd0):(4'd4))));
  localparam [3:0] p12 = (~^((3'sd0)?(&(^(2'd0))):(~(~|(-2'sd0)))));
  localparam [4:0] p13 = {1{(!(|(~({2{(4'd9)}}!==((-2'sd0)===(2'd3))))))}};
  localparam [5:0] p14 = (((4'd2 * (4'd0))&((5'sd13)!==(4'd2)))^{2{((2'd3)||(3'd7))}});
  localparam signed [3:0] p15 = (((~(5'd17))>=(2'd3))+(4'sd1));
  localparam signed [4:0] p16 = {3{(2'd3)}};
  localparam signed [5:0] p17 = {2{{3{(2'd1)}}}};

  assign y0 = (~&(a1<=a3));
  assign y1 = ((~|(-$unsigned($signed($signed((~^(+($signed((~^($unsigned(a2)))))))))))));
  assign y2 = (({(b0>>>p14)}^({p0}+(5'd2 * b1)))+(({a5}>>>(p8<<<p14))&&{p10,p16,p5}));
  assign y3 = ((-((&a4)?(p17<<p4):(+p15)))?(5'sd14):(~^(~(p4?b2:p6))));
  assign y4 = $signed((p0>p0));
  assign y5 = ({4{{3{p8}}}}&&(((b2|a1)!=={1{a4}})));
  assign y6 = (^{{a2,b5},(a2!==b3),(3'd7)});
  assign y7 = (&((&(~^a5))||(p16|p4)));
  assign y8 = ((-2'sd1)%p15);
  assign y9 = ((((a5<a2)^(p10>p5))<<<((a3===a4)-(a3<b0)))>>(^{{a1,p9},(~|(^b2)),(b4^p2)}));
  assign y10 = ((5'sd10)?{p9,p11}:{p7,p10,b2});
  assign y11 = (&{4{p9}});
  assign y12 = ((b0?p1:b2)+(p1<=a2));
  assign y13 = (p5==p12);
  assign y14 = ((2'sd1)?{2{p2}}:(a4!==a3));
  assign y15 = (~|$signed({{2{(p16&b5)}},((b5===b0)>(|$unsigned(p9))),{(+(&$signed((|b1))))}}));
  assign y16 = (({(a4<<p14),(b1!==a2)}|(4'd9))^(-2'sd1));
  assign y17 = {(b4),{p8,p10},(p6||a1)};
endmodule
