module expression_00567(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd5)<=(4'd0));
  localparam [4:0] p1 = ((4'd2 * {3{(3'd7)}})^{2{({(4'd2),(3'd2)}!={(-4'sd3)})}});
  localparam [5:0] p2 = (-{4{(3'd2)}});
  localparam signed [3:0] p3 = ((+(3'sd0))==((4'sd1)<<<(3'd6)));
  localparam signed [4:0] p4 = ((2'sd1)>>>(5'sd11));
  localparam signed [5:0] p5 = (((2'sd1)==(5'd22))>>(~&(-(3'd1))));
  localparam [3:0] p6 = (((2'd1)?(-4'sd6):(3'd1))%(5'sd13));
  localparam [4:0] p7 = ((2'd2)^((2'd2)|(3'sd2)));
  localparam [5:0] p8 = ({(3'd0),(-5'sd11),(4'd10)}?((3'sd3)|(5'd1)):{(5'sd5),(3'sd0),(2'sd0)});
  localparam signed [3:0] p9 = ({(-3'sd2),(2'd1),(3'd6)}!==(((5'd0)>>>(-5'sd6))<{(3'd6)}));
  localparam signed [4:0] p10 = (2'sd1);
  localparam signed [5:0] p11 = ((5'd14)?(~|(&((5'd15)?(-2'sd0):(5'd26)))):{(3'd4),(5'sd12),(2'd0)});
  localparam [3:0] p12 = {((+(4'sd1))?(!(4'sd0)):{(-4'sd4),(-4'sd0),(-2'sd0)})};
  localparam [4:0] p13 = (((~|{(3'd3)})^~((4'd14)>>(2'd3)))!==(6'd2 * {((5'd14)<<(2'd0))}));
  localparam [5:0] p14 = {{{{(4'sd4),(5'sd0)},{(2'd1)}}}};
  localparam signed [3:0] p15 = ((2'd1)|(-5'sd9));
  localparam signed [4:0] p16 = ((3'sd3)-(3'sd0));
  localparam signed [5:0] p17 = (-5'sd10);

  assign y0 = (~^((5'sd1)>=(~&(p1||p4))));
  assign y1 = {1{({4{{1{p2}}}}>={1{({3{b4}}<<(a5==b4))}})}};
  assign y2 = ((($signed($unsigned($signed(p7)))^~((p8&p11)<<(p1))))<($signed(((a1==a2)+(a1===a2)))!==(($unsigned(a3)-$unsigned(b1)))));
  assign y3 = (2'd2);
  assign y4 = (-{4{(!b1)}});
  assign y5 = ((~|b0)?(^p13):(-a2));
  assign y6 = ((3'd2)>{a2,p1,p14});
  assign y7 = (!((-3'sd3)^(~(^(+a5)))));
  assign y8 = {3{{2{{1{a2}}}}}};
  assign y9 = {(!((p3&&p13))),((&b1)+{a2})};
  assign y10 = {2{{4{a4}}}};
  assign y11 = ({(p11>=p16),(p2?p8:p14),(-p1)}?((p1)>>>(p10&&p11)):((-p14)|(2'sd1)));
  assign y12 = ($unsigned((&$signed((2'd1))))>>(-(((a0-a1))<<<((~&p12)+(~|p10)))));
  assign y13 = (^(~|((b5>>a2)<<<(a4>>p0))));
  assign y14 = {(5'd16),(((a0-p4)<<<{p5})&&((3'd7)-(-2'sd0)))};
  assign y15 = (-2'sd0);
  assign y16 = (((+(+(b4&p3)))+({b1,p5,b3}?(p12-p17):(a0?p5:p6)))^~((&(p13|p8))?(^(+p16)):{(a5?a4:a0)}));
  assign y17 = {{2{(p17?p10:p15)}},($unsigned((p7^p16))+(p14>=p9))};
endmodule
