module expression_00286(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^((5'sd14)?(3'd2):(-4'sd0)));
  localparam [4:0] p1 = (~&((-3'sd1)>=(&(2'd2))));
  localparam [5:0] p2 = (4'd14);
  localparam signed [3:0] p3 = (~{2{{4{(5'd27)}}}});
  localparam signed [4:0] p4 = (~(5'd14));
  localparam signed [5:0] p5 = (~^(((4'sd4)>>>(-2'sd0))===((-4'sd7)!=(-5'sd0))));
  localparam [3:0] p6 = (-4'sd3);
  localparam [4:0] p7 = ((-(+(3'd2)))?((3'd3)?(5'sd2):(2'd2)):((-4'sd2)?(2'd3):(-5'sd13)));
  localparam [5:0] p8 = (^(5'd27));
  localparam signed [3:0] p9 = {1{(-2'sd1)}};
  localparam signed [4:0] p10 = ({1{(((-5'sd13)!==(3'sd2))^{3{(4'sd5)}})}}<<<{2{(~(-3'sd2))}});
  localparam signed [5:0] p11 = ((4'd10)>>{3{(2'd2)}});
  localparam [3:0] p12 = (({1{(~(3'd4))}}<<<(^{1{(5'sd10)}}))>>(((5'sd8)<=(2'd0))?((2'sd0)<=(2'd1)):((5'd16)&&(-2'sd1))));
  localparam [4:0] p13 = ((5'd0)?((4'sd4)&&(2'd0)):(-4'sd2));
  localparam [5:0] p14 = (~((((2'd0)<(5'd27))!==((4'sd4)?(4'd9):(-3'sd1)))&&{((-3'sd1)?(5'd18):(-5'sd0)),((5'sd5)?(-3'sd2):(3'sd1))}));
  localparam signed [3:0] p15 = ({3{((2'd3)?(2'd3):(5'sd3))}}>=((~(-3'sd0))|((5'd3)<<(4'sd0))));
  localparam signed [4:0] p16 = ((-5'sd2)^~(~|(5'sd4)));
  localparam signed [5:0] p17 = (((4'd15)^~(-4'sd7))>>>(2'sd1));

  assign y0 = (((p17?p15:p9)|(4'd2 * a2))?(~{2{(a3>>p6)}}):((!a4)===(^b3)));
  assign y1 = {4{(5'sd7)}};
  assign y2 = (p4?b3:a1);
  assign y3 = {3{({3{b0}}!=$unsigned(p9))}};
  assign y4 = $unsigned($unsigned({3{(5'd28)}}));
  assign y5 = $unsigned($signed((((p8-p17))<<<(~|(p6/p4)))));
  assign y6 = (5'd2 * $unsigned((4'd0)));
  assign y7 = {p0,p3,p12};
  assign y8 = ((p1&&p7)<<<(p17||p7));
  assign y9 = ((p7||p11)|(|p16));
  assign y10 = {2{(2'sd0)}};
  assign y11 = ((&(6'd2 * (~|{4{b1}})))?((p2?a2:a1)&&(b3^p16)):$unsigned((~&(~(-(a1>>p6))))));
  assign y12 = {4{{{3{b5}},{b5}}}};
  assign y13 = (((&b1)<(^a3))!==(~(b3>b5)));
  assign y14 = (&(!(^$unsigned({4{$signed({4{b2}})}}))));
  assign y15 = (~^(({3{$unsigned(p6)}}?((|(!p11))^~{2{p3}}):({3{a1}}?$signed(p4):(a1^~p1)))));
  assign y16 = ({a3,b0,b3}+{a1});
  assign y17 = (-2'sd1);
endmodule
