module expression_00003(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-{2{{4{(2'd3)}}}});
  localparam [4:0] p1 = (2'sd0);
  localparam [5:0] p2 = {((5'd26)?(3'd4):(2'd1)),((3'sd3)?(3'd2):(3'd4)),((2'd3)?(-4'sd6):(4'd6))};
  localparam signed [3:0] p3 = (~&(((3'sd3)?(3'd7):(2'sd1))?({(3'd2)}^~((-2'sd1)|(-5'sd13))):((4'd2 * (5'd6))=={(4'd15)})));
  localparam signed [4:0] p4 = (~^{2{((^{2{(5'sd9)}})==(5'd26))}});
  localparam signed [5:0] p5 = {{2{{(4'd11),(-3'sd1)}}}};
  localparam [3:0] p6 = ((((3'sd0)&&(2'd1))*((5'sd5)===(-5'sd7)))<<(((4'sd4)>>(2'sd0))/(-3'sd3)));
  localparam [4:0] p7 = ((5'd9)|(4'sd2));
  localparam [5:0] p8 = (|((2'sd1)?{1{(3'd5)}}:(-(5'd20))));
  localparam signed [3:0] p9 = {1{(+{4{(4'd1)}})}};
  localparam signed [4:0] p10 = (~|(({4{(4'd4)}}?(+(5'd22)):(~(5'sd12)))?(^(~&{2{(4'sd3)}})):(((4'd10)?(3'sd1):(5'd12))?(~&(3'sd1)):((-5'sd9)?(4'd7):(5'd30)))));
  localparam signed [5:0] p11 = {(-3'sd2),(5'sd2),(-5'sd14)};
  localparam [3:0] p12 = {4{(2'd0)}};
  localparam [4:0] p13 = (+(~&({2{{(-5'sd8),(2'd2)}}}-({(2'd2),(5'd2),(3'sd1)}<<{3{(4'd4)}}))));
  localparam [5:0] p14 = {({1{((5'd7)>>(-4'sd5))}}?(6'd2 * (5'd16)):{(5'd28),(4'd11),(2'sd0)})};
  localparam signed [3:0] p15 = ((((4'sd0)^~(3'd3))>((3'd7)+(-3'sd2)))&(&(((5'sd0)===(3'd5))>>>(~(3'd0)))));
  localparam signed [4:0] p16 = (-2'sd1);
  localparam signed [5:0] p17 = (&(-(-((~(^{(+(4'd15)),{(-5'sd11),(2'd0),(2'sd1)}}))||(!(((4'sd6)>(5'sd5))<=(2'sd1)))))));

  assign y0 = ({1{(2'd3)}}>>>(b0^a1));
  assign y1 = (~&{((~|(a5>b5))!==(b0>>>b4)),(~&(5'd2 * (p2>=b2))),((^(4'd2 * p1))>>>(b1==b3))});
  assign y2 = (({a1}^~{b5,b0})===((|b1)==={a4}));
  assign y3 = (((p5^~p12)||($unsigned(b4)))?(((p3?p17:p3)?(p11<<p16):(p3>p7))):($signed(a4)?(p16>>a5):(b0?p3:a0)));
  assign y4 = ((p6?p9:p14)?(p7?p3:p10):(p6<<<p9));
  assign y5 = ({{2{b0}}}!=={3{b1}});
  assign y6 = (-(-(+{((+(!(-p9)))^{(4'd2 * p13),{p1,p6}}),(((!p17)+(!a4))|(~&{a2,p13}))})));
  assign y7 = (!{3{(p12&&a4)}});
  assign y8 = (&({3{b4}}?(~(p0?a2:p17)):(-{2{p15}})));
  assign y9 = (a4&&p16);
  assign y10 = ({(p12^p17),(p5<<a5),(~&(p8!=p5))}>=(^(-{{(~b1),{a5,a1}},((|a4)<=(p12==p12))})));
  assign y11 = ((a1&p12)?(p6^~p6):(b0!=p8));
  assign y12 = (^(4'sd7));
  assign y13 = $unsigned(($signed(b5)));
  assign y14 = (p0?p13:p3);
  assign y15 = {{(~|(~&b0)),{p3,p15}},(~&{2{{3{p3}}}})};
  assign y16 = (~(5'd18));
  assign y17 = {{(~&{{2{p8}},(~&p4),(~^p6)}),({1{(p16!=p15)}}!=(b0===b3)),({1{(p17+p5)}}<={2{p6}})}};
endmodule
