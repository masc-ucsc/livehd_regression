module expression_00109(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(&(4'd9)),(-3'sd1)};
  localparam [4:0] p1 = {4{((3'd3)?(3'd2):(-2'sd0))}};
  localparam [5:0] p2 = ((((4'd11)==(2'd3))/(4'd10))>>(((-3'sd3)?(-3'sd2):(-3'sd0))<<(-((-2'sd0)?(3'sd3):(5'd11)))));
  localparam signed [3:0] p3 = {(2'sd0),(5'd11),(5'd17)};
  localparam signed [4:0] p4 = (^((~(4'd13))?{4{(-2'sd0)}}:((2'sd1)?(5'sd9):(4'd14))));
  localparam signed [5:0] p5 = (^{2{(2'd0)}});
  localparam [3:0] p6 = ({3{(-3'sd3)}}>=((5'd5)^(-3'sd0)));
  localparam [4:0] p7 = {(3'd4),(5'd9),(2'd1)};
  localparam [5:0] p8 = (({2{((3'sd0)==(2'd1))}}<<<(((3'sd2)<<<(2'd3))<<<((4'd5)===(4'sd2))))&&(^(&(((4'sd5)>(-4'sd0))-{1{((4'd5)^~(-2'sd0))}}))));
  localparam signed [3:0] p9 = (^((~|(~((+(4'd6))<<(~^(-3'sd3)))))<=(3'sd3)));
  localparam signed [4:0] p10 = ((-3'sd0)^~(5'd8));
  localparam signed [5:0] p11 = (((3'sd3)>>>(4'd14))?((3'sd0)?(4'sd5):(-2'sd0)):((-2'sd0)?(4'd14):(5'sd11)));
  localparam [3:0] p12 = (|(&(&{(&{(3'd4)}),(+(~^(-4'sd3))),(6'd2 * (3'd2))})));
  localparam [4:0] p13 = (4'sd7);
  localparam [5:0] p14 = ((^(&(2'd2)))==={((4'd11)-(-4'sd6))});
  localparam signed [3:0] p15 = ((3'sd3)?(5'sd4):(3'sd3));
  localparam signed [4:0] p16 = {(-{((~^(5'd19))?((3'd5)?(2'sd1):(4'd4)):{(2'd1)})})};
  localparam signed [5:0] p17 = (({4{(2'd1)}}||(5'd28))>=(4'd15));

  assign y0 = (+(-(~&(!(~|(!(b4<<<p15)))))));
  assign y1 = {4{(6'd2 * (a2&&a2))}};
  assign y2 = (((&p16)>(~&b3))<=({p4}||(a2-b0)));
  assign y3 = $unsigned(((((b1)-(5'd2 * p13))|$signed((a0>>>p8)))+($unsigned($signed($signed(p12)))<<<((a5&&b5)===(b4&&b0)))));
  assign y4 = ((~|(p0&b3))>>>((a2||a4)<(^b3)));
  assign y5 = ((((b3<<<a2)<=(p16*p6))>=((b1/a5)!=(p4^a0)))^(((p5&&b0)&(b1%p13))>>>((p0^b3)||(b1===a0))));
  assign y6 = {1{$signed((-2'sd0))}};
  assign y7 = (!(+({a5,b1}<<<{a0,a3})));
  assign y8 = {((~&(b2>>p0))||(^(p14||p3))),{({a2,p0,a2}<<{4{p8}}),{(+(4'd11))}}};
  assign y9 = (+(((&b0)?{3{b1}}:(a3?b3:a3))?({4{b0}}|(a0?a4:b2)):({3{a4}}<<<(a1&b2))));
  assign y10 = {4{a0}};
  assign y11 = (~&(p17>>b2));
  assign y12 = $signed((4'sd3));
  assign y13 = ($unsigned(((b3&a3)<<$signed(p1))));
  assign y14 = ({{p1,p2},{p7,p17,p3},(p12^p10)}&&((|p14)?(~|p8):(2'sd0)));
  assign y15 = (~^(((~|(a3<<a2))<<<(-3'sd3))^~(~^(3'd1))));
  assign y16 = (|{a1,b2,p6});
  assign y17 = (((a0+a1)|(b2<<<a3))&&((~&p12)||{4{p9}}));
endmodule
