module expression_00144(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({{(-5'sd14),(5'sd3),(-2'sd0)},((-5'sd11)|(3'd3)),((5'd10)|(5'sd0))}?{{(3'd4),(-2'sd0)},((4'd0)>>>(4'sd5)),(5'd2 * (3'd3))}:(((3'd1)<<<(-2'sd1))|((4'd13)?(3'd3):(5'sd5))));
  localparam [4:0] p1 = {1{((4'sd5)^~(-2'sd1))}};
  localparam [5:0] p2 = (&{(4'd2 * ((5'd17)^(2'd1)))});
  localparam signed [3:0] p3 = {3{((5'sd12)-(2'd2))}};
  localparam signed [4:0] p4 = (+(^(~^(5'd7))));
  localparam signed [5:0] p5 = {{(3'sd2),{(-5'sd1)}},{{(3'd4)},{(-5'sd15)}},{{(5'd9),(5'd3),(3'd6)},(2'd3)}};
  localparam [3:0] p6 = (-(-(4'sd4)));
  localparam [4:0] p7 = {1{(2'sd1)}};
  localparam [5:0] p8 = ((~&(^(((-5'sd1)*(5'd17))>>(~(2'd0)))))===((~|(~&(5'd18)))>=((3'd1)?(-5'sd14):(4'sd0))));
  localparam signed [3:0] p9 = (-4'sd4);
  localparam signed [4:0] p10 = (2'sd1);
  localparam signed [5:0] p11 = (-5'sd2);
  localparam [3:0] p12 = ({1{{3{(4'd15)}}}}!=(((3'd2)||(-3'sd0))>>{4{(5'd0)}}));
  localparam [4:0] p13 = {(3'd5),(5'd3)};
  localparam [5:0] p14 = (4'sd7);
  localparam signed [3:0] p15 = ((5'sd0)!=(5'sd7));
  localparam signed [4:0] p16 = {(-4'sd5),(5'd5)};
  localparam signed [5:0] p17 = ((((-5'sd8)^~(-2'sd0))<{((-3'sd0)!==(3'd1))})!={((4'sd7)!=(4'sd0)),((2'sd0)<<(2'd3)),(~(5'd18))});

  assign y0 = (-(!p4));
  assign y1 = ((p11?b5:a0));
  assign y2 = {2{(-3'sd1)}};
  assign y3 = (5'd4);
  assign y4 = (3'sd1);
  assign y5 = {4{(a1===a0)}};
  assign y6 = ((~^$signed((-2'sd1))));
  assign y7 = ((p8==p4)?(p7?p5:p3):(a5!==b3));
  assign y8 = (~|(((a2&&p11)==(a1<a0))?((a0?b1:b1)?(b2&&b3):(-2'sd1)):(^((+b3)<=(~|a0)))));
  assign y9 = (&(((^(($unsigned(p1)!=(!b0)))))+(~(+(|(~{3{b4}}))))));
  assign y10 = (5'd2 * (4'd11));
  assign y11 = (~^(3'd3));
  assign y12 = (4'd2 * (p7+b1));
  assign y13 = (($unsigned(a1)?$signed(p1):{1{b3}})||((5'd14)));
  assign y14 = ((b5|b4)%b4);
  assign y15 = (4'd11);
  assign y16 = (~(((a3!==b4)||(a2^b0))));
  assign y17 = (~&(-5'sd9));
endmodule
