module expression_00998(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd0);
  localparam [4:0] p1 = ((3'd7)?(3'sd0):(-2'sd1));
  localparam [5:0] p2 = ((-3'sd0)>=(((5'd2)<<(5'sd11))<((3'd3)^~(-3'sd3))));
  localparam signed [3:0] p3 = (~^((~^({4{(5'sd10)}}>>>{4{(4'd2)}}))<<(~{2{(&(3'sd3))}})));
  localparam signed [4:0] p4 = ((((3'sd0)||(2'd1))==={(2'd2)})<{{(3'd5)},((2'd1)|(4'sd1)),{(-4'sd4),(3'sd2)}});
  localparam signed [5:0] p5 = (-4'sd5);
  localparam [3:0] p6 = (^{3{(5'd25)}});
  localparam [4:0] p7 = (({4{(4'sd1)}}>((-2'sd0)+(-2'sd1)))<={(5'd30),(3'd2),(4'd8)});
  localparam [5:0] p8 = {2{(5'sd5)}};
  localparam signed [3:0] p9 = ((((4'd0)*(3'sd1))?((3'd4)===(-4'sd7)):((-5'sd2)<<(-5'sd8)))^(((2'd0)?(2'd0):(3'd5))%(4'sd1)));
  localparam signed [4:0] p10 = {1{(({(4'd1),(5'd9)}==={2{(2'd1)}})!==((6'd2 * (5'd23))>{4{(-4'sd2)}}))}};
  localparam signed [5:0] p11 = {2{({2{(2'sd1)}}<(-(-4'sd5)))}};
  localparam [3:0] p12 = ((4'd11)>(2'd0));
  localparam [4:0] p13 = (6'd2 * ((3'd0)%(4'd4)));
  localparam [5:0] p14 = ({{(-5'sd13),(2'd2),(2'd2)}}?({(3'sd3),(4'sd5),(3'd1)}?{3{(-4'sd6)}}:((5'd4)?(-5'sd4):(5'd27))):{3{{3{(5'd24)}}}});
  localparam signed [3:0] p15 = (((5'd14)?(5'sd15):(4'sd7))<<<(!((3'd1)?(3'sd3):(5'd17))));
  localparam signed [4:0] p16 = (|(3'd5));
  localparam signed [5:0] p17 = (~&(4'd9));

  assign y0 = $unsigned(a2);
  assign y1 = ((4'sd6)?(p13):(p10?p13:p9));
  assign y2 = (2'd0);
  assign y3 = {3{(+((b1?p2:a5)?(p1||a5):(a2!==b3)))}};
  assign y4 = (^(((~|{3{{2{p17}}}})||((-2'sd1)+{a0,p1}))));
  assign y5 = (^{1{(^{(~&{1{p7}}),(p4<<b0),(p11<<<b1)})}});
  assign y6 = $signed({{p9,a3,p3}});
  assign y7 = ((4'd2 * (b1^b0)));
  assign y8 = (|((2'sd1)||(~^(!(p3?b4:b3)))));
  assign y9 = (!(~^((p16?a3:p8)?(a3&p1):(a2&&p16))));
  assign y10 = {(p4<<p0),(p6-p3),(p10?b5:p7)};
  assign y11 = $unsigned(((p5?a0:b2)?(|(-(p9))):((p4?p9:p17)==(p4==p7))));
  assign y12 = ($signed({1{p14}})!=(a4?a3:a3));
  assign y13 = (((~&p2)?{1{p17}}:(+p9))^~(~((~^p10)?(b5?p16:b4):(a2?p6:b3))));
  assign y14 = ({((|{(b3^p12)})?(({3{p3}})):(|(~^(~&$unsigned(p15)))))});
  assign y15 = ((a3<<<a5)>(^a4));
  assign y16 = {b2,p12,p8};
  assign y17 = $signed(({4{(|(p10&&p11))}}));
endmodule
