module expression_00319(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(^(3'd5))};
  localparam [4:0] p1 = {(!(3'd4))};
  localparam [5:0] p2 = ((~^(((2'd1)!=(2'd3))!==((3'd7)>=(4'd3))))<<<((+((5'd1)<<<(-2'sd1)))%(5'sd5)));
  localparam signed [3:0] p3 = {{(2'd3),(2'd1),(2'd2)},{4{(4'd2)}}};
  localparam signed [4:0] p4 = ({(-4'sd6)}-(~&({(3'sd2),(-3'sd1)}^{(2'd0),(-2'sd1)})));
  localparam signed [5:0] p5 = {{(2'd2),(4'sd4),(4'd1)},{1{((4'd6)|(4'sd4))}},((4'd11)?(-4'sd3):(-3'sd0))};
  localparam [3:0] p6 = ({(|(-5'sd9)),(^(3'd2)),{(-4'sd4)}}&&(-((-2'sd0)<((-4'sd1)&&(3'd0)))));
  localparam [4:0] p7 = ((!((&(5'd21))?((2'd1)?(2'd1):(3'd0)):{(-4'sd0)}))^~(((-5'sd9)?(4'd1):(5'd12))!=(5'd6)));
  localparam [5:0] p8 = {1{((-3'sd2)&(4'd10))}};
  localparam signed [3:0] p9 = (3'd4);
  localparam signed [4:0] p10 = (((2'd1)-(4'd12))?((2'sd0)===(3'd3)):(4'd8));
  localparam signed [5:0] p11 = (!((~((|(5'd11))<((4'd5)^(3'd1))))+(^(~^((5'sd12)^~(2'd2))))));
  localparam [3:0] p12 = (~^{2{{(~^((5'd15)==(-2'sd0))),((5'd30)&&(5'd23))}}});
  localparam [4:0] p13 = (((-4'sd5)<=(5'd23))!=((-5'sd6)>>(4'd12)));
  localparam [5:0] p14 = (5'd2 * ((2'd1)||(5'd19)));
  localparam signed [3:0] p15 = (5'd12);
  localparam signed [4:0] p16 = (((5'sd8)&(5'd20))?((2'sd1)?(5'sd7):(2'd0)):{((4'sd0)<<(4'd6))});
  localparam signed [5:0] p17 = ((5'd22)^((2'd2)^(2'd2)));

  assign y0 = ({2{p0}}?(p7!=p2):{4{a0}});
  assign y1 = {3{(~&{b2})}};
  assign y2 = ((5'd2 * (p8||p14))^~(((p4<<p6)<=(p14>=p3))^~((p8>=p0)&&(|a5))));
  assign y3 = ({((b1?b2:b0)===(a5?a5:b1))}-((p17-p10)!={p1,p14,p8}));
  assign y4 = ((~&(p9?p4:p17))?(!$signed((-(!p16)))):((|a5)!==$signed(b1)));
  assign y5 = $signed({(a0-p11),(a3==a0),(p13)});
  assign y6 = (((6'd2 * (p6/a0)))^~(((a3|a2)|$unsigned(a0))==(~(!(b2===b2)))));
  assign y7 = (((4'd2 * a2)+(a5!=b5))<=((b1!=a0)=={a5}));
  assign y8 = ({(~^(3'd0)),(&(&a0)),(2'd1)}==={({(~|(&b3))}<<(b5?b4:a1))});
  assign y9 = ({4{{3{p5}}}}<<{{{a5,a1,p5},(p0^~p17)}});
  assign y10 = {{($signed(a3)?{a3,a2}:(a3+p16)),({p4}>>>(b4>>>a5)),{{a2,a2,a5},(|a0),{b3,a1}}}};
  assign y11 = $unsigned(((b3?a1:p14)<$unsigned(p8)));
  assign y12 = ((2'sd0)%p4);
  assign y13 = {((p8||p8)?{{p10}}:(p8||p16)),(4'd13)};
  assign y14 = {a0,b4,b4};
  assign y15 = {(-2'sd0),({b1,a1}<=(~&p14))};
  assign y16 = {($signed(((b4<<a3)===(b5&b0)))),(^{{1{{3{p8}}}},(!(b1&a0)),{3{a2}}})};
  assign y17 = {1{(2'd1)}};
endmodule
