module expression_00642(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd0)?(-4'sd4):(-3'sd1))||((2'd0)?(4'd5):(5'd7)));
  localparam [4:0] p1 = (((((2'sd0)?(4'd8):(4'd13))>>>((3'sd2)^(5'd21)))||(((5'sd5)^~(-3'sd1))>((2'd0)?(3'd4):(-3'sd3))))===(+(((2'sd0)^~(2'd1))^~((2'sd1)<<<(3'd6)))));
  localparam [5:0] p2 = (~&{(4'd2 * (5'd15)),(~&{(2'd2)})});
  localparam signed [3:0] p3 = (4'd2 * ((2'd1)-(3'd4)));
  localparam signed [4:0] p4 = ((3'sd0)?((4'sd4)?(5'sd8):(5'd8)):(~((2'sd1)?(5'sd13):(4'd8))));
  localparam signed [5:0] p5 = (((!((3'sd2)>>(5'd18)))!=={(2'd0),(5'd19)})+({3{(-4'sd7)}}<<<((4'd2)&&(3'sd0))));
  localparam [3:0] p6 = (&(~^(~(-(~|(~&(|(3'd3))))))));
  localparam [4:0] p7 = ((5'd5)<=(4'd10));
  localparam [5:0] p8 = ({(4'd13),(-5'sd13),(4'd7)}<<<(~^((5'd27)<(4'sd3))));
  localparam signed [3:0] p9 = (((-2'sd0)?((5'd6)?(4'd2):(4'sd7)):(4'd13))>>>(((3'd5)?(4'd8):(-3'sd3))?(2'sd1):((-4'sd3)?(2'd3):(4'd2))));
  localparam signed [4:0] p10 = ({1{(((-3'sd1)?(3'd2):(2'sd1))!==(^(5'd7)))}}!={1{(-2'sd1)}});
  localparam signed [5:0] p11 = (-3'sd2);
  localparam [3:0] p12 = (((-4'sd3)<<<(2'sd1))!==((4'sd3)<=(4'd8)));
  localparam [4:0] p13 = (4'd0);
  localparam [5:0] p14 = (~^((^(&((4'sd0)!=(!(4'd2)))))^~((~^(2'sd1))+((5'sd11)*(2'd0)))));
  localparam signed [3:0] p15 = ({4{(5'sd5)}}?(~&{3{(3'sd2)}}):(!((3'sd0)>>(-5'sd6))));
  localparam signed [4:0] p16 = (!(2'sd0));
  localparam signed [5:0] p17 = ((((5'd18)/(5'sd15))/(5'd12))?((-3'sd3)|((-2'sd0)%(2'd3))):(-2'sd1));

  assign y0 = (3'd6);
  assign y1 = (!$unsigned((3'sd2)));
  assign y2 = (2'd3);
  assign y3 = ((+((b5<=a2)?(b5>=p8):(^b1)))?((-(b4?a0:a4))+(a4==a5)):((b3?a0:b2)?(~^a5):(a2?a3:a2)));
  assign y4 = (((3'd1)^((5'd24)+(a4&&b5)))+(2'd2));
  assign y5 = (2'd0);
  assign y6 = (~|(4'sd1));
  assign y7 = ((~(&((~(p7>>p12))+(+(4'd9)))))^((-(p12|p17))==(-(-3'sd2))));
  assign y8 = $signed((~^(((p6)<<(p16&p15))>>>(~{2{a3}}))));
  assign y9 = (-((5'd1)?(4'd2 * (3'd6)):((a1?a1:a1)&(p17^~b4))));
  assign y10 = {((b0>a0)^~(b3>>a3)),($signed({p10,b4,b3})<<<(p2?a2:p7)),$signed(($unsigned((b0|b0))!=(b3?p13:a2)))};
  assign y11 = $unsigned(({((p7)^(p4<b5)),({b4,a5}!=(b0||b4))}|(((p2<=p7)>(p3>>p7))-(+{p11,p9,p2}))));
  assign y12 = (p8?b5:p5);
  assign y13 = (4'd2);
  assign y14 = {2{$unsigned((b0?a1:b5))}};
  assign y15 = ((a0!==a0)&(b0?p12:p5));
  assign y16 = ((2'sd1)>=(-2'sd0));
  assign y17 = (({4{p3}}||((b3!=p13)&(a4?p2:p6)))&(((p12<p4)<<(p15?p15:p4))<(a1?p1:p15)));
endmodule
