module expression_00264(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{{(3'sd2),(3'sd2),(5'd29)},{(5'd9),(5'd9)}}};
  localparam [4:0] p1 = (({4{(5'd5)}}!==((-2'sd1)?(4'sd1):(4'd3)))<<{1{(((5'sd4)?(5'sd1):(5'sd6))&&((5'sd13)?(2'sd0):(2'd0)))}});
  localparam [5:0] p2 = {(2'sd0)};
  localparam signed [3:0] p3 = ((3'd6)?(2'sd0):(3'd6));
  localparam signed [4:0] p4 = {(~^{{1{{2{{3{(2'd2)}}}}}}})};
  localparam signed [5:0] p5 = ((3'd1)||(5'd30));
  localparam [3:0] p6 = (~^(5'd18));
  localparam [4:0] p7 = ((-5'sd2)&&(2'd1));
  localparam [5:0] p8 = {(((-5'sd1)>>(-2'sd0))&((4'sd3)?(2'sd1):(4'd11))),((5'd22)?(5'sd0):(3'd4)),{((5'd21)>>>(2'd2))}};
  localparam signed [3:0] p9 = ((-2'sd0)^~(((3'd5)?(-5'sd8):(-4'sd2))!=(3'sd0)));
  localparam signed [4:0] p10 = {(2'd1)};
  localparam signed [5:0] p11 = (-((~(~|(~&{3{(-2'sd0)}})))<(((-2'sd0)?(2'd1):(3'd7))?((4'd3)==(-2'sd0)):(-(3'd3)))));
  localparam [3:0] p12 = {{(2'd2),{(4'd10),(3'd1),(4'sd7)}},(4'd0)};
  localparam [4:0] p13 = (((-3'sd3)?((4'sd7)-(5'd31)):(5'd12))>=((5'd7)+(-4'sd2)));
  localparam [5:0] p14 = ((2'sd1)^(3'd1));
  localparam signed [3:0] p15 = (~&{2{({(-2'sd1),(4'd15)}&{3{(-3'sd0)}})}});
  localparam signed [4:0] p16 = {(|(~(-4'sd4))),((4'sd5)|(4'd13)),(!{(2'd0),(4'd2),(-2'sd1)})};
  localparam signed [5:0] p17 = (-5'sd2);

  assign y0 = (((b2!==b4)+(|a3))+($unsigned(p5)>>>(-2'sd0)));
  assign y1 = {((^p3)?(+p10):{p3,p16,p7}),(+((&a4)==={a4}))};
  assign y2 = (5'sd4);
  assign y3 = (((-{(((a2===b5))||(a0&&b1))}))==(^(&((p3?p6:b1)>>($unsigned(a4)<=(+a2))))));
  assign y4 = {4{$signed((p3))}};
  assign y5 = {2{$unsigned($unsigned((((b5?a3:a5)<<(|a0))||(4'd2 * (~&a1)))))}};
  assign y6 = (^(-(+(+{b5}))));
  assign y7 = ({2{(p13?p10:p12)}}?((~|(5'd22))>>(p2?p6:p6)):((p5^p1)&(p11^~p11)));
  assign y8 = (p7<<<p17);
  assign y9 = (-5'sd5);
  assign y10 = (~|(((~(&a5))<<(a4^~b2))!=={{(a4),(a0^~a5),(a1>>b0)}}));
  assign y11 = ((~((6'd2 * a2)|(a2<=p16)))>=((p17<<b0)*(b5+p0)));
  assign y12 = (5'sd6);
  assign y13 = (~(-(|(~^(~|(|(p14>>>p0)))))));
  assign y14 = {4{(~&{p16,p9,p12})}};
  assign y15 = ((6'd2 * (b0===b2))!==((a4?a4:a3)&(|b1)));
  assign y16 = ((-2'sd1)&(6'd2 * p1));
  assign y17 = {4{$unsigned(((a1<p4)))}};
endmodule
