module expression_00464(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({1{(5'd24)}}>>{4{(4'sd2)}})!==(-4'sd1));
  localparam [4:0] p1 = ((5'd2 * (5'd11))^~{2{(4'd15)}});
  localparam [5:0] p2 = (|(~^{(!(-3'sd2)),(^(4'sd4))}));
  localparam signed [3:0] p3 = (((4'd14)*(4'sd4))^((-3'sd1)>=(5'sd12)));
  localparam signed [4:0] p4 = {(^(3'd7)),(2'd3)};
  localparam signed [5:0] p5 = (5'd2 * ((4'd4)&&(4'd12)));
  localparam [3:0] p6 = (~|{1{(((5'd19)<(5'd22))||(-(5'd31)))}});
  localparam [4:0] p7 = ({4{(2'd1)}}?{(2'd3),(5'd6),(2'd1)}:{((5'd7)?(-2'sd0):(-2'sd1)),((4'd14)|(4'd13))});
  localparam [5:0] p8 = ({((-3'sd0)^(-5'sd9)),((5'd23)?(4'd9):(-4'sd3)),{1{((5'd10)?(5'd30):(2'sd1))}}}!=({(5'd2 * (2'd2))}^(~&((4'd3)?(4'd3):(5'sd13)))));
  localparam signed [3:0] p9 = (~&(-5'sd0));
  localparam signed [4:0] p10 = (~|(~(^(-(&{(+(^{{(2'd1),(2'd3),(2'd2)},{(5'd30)},{(5'sd12)}}))})))));
  localparam signed [5:0] p11 = (!(^(-4'sd0)));
  localparam [3:0] p12 = (~{1{(2'd2)}});
  localparam [4:0] p13 = (4'd2 * ((5'd29)?(3'd1):(5'd1)));
  localparam [5:0] p14 = (3'd6);
  localparam signed [3:0] p15 = (({2{(-5'sd11)}}&((-4'sd7)-(5'd0)))<<<{2{{2{(2'd0)}}}});
  localparam signed [4:0] p16 = (~|{(~&(~|(5'd2))),(2'd2),((5'sd15)+(-4'sd0))});
  localparam signed [5:0] p17 = (2'sd1);

  assign y0 = (~(&((+(~&(p12>a5)))>{{2{(|a2)}}})));
  assign y1 = (~^(~^(5'd15)));
  assign y2 = (-(+((!((~^(a1?p11:a2))>>>(p1||p3)))<<(|({4{p3}}<={p1,b1})))));
  assign y3 = (-(^{2{(-(4'sd4))}}));
  assign y4 = ($unsigned((4'd2 * {p14,a0,b0}))||{{(a5<b2),(b0===b2),$unsigned(p12)}});
  assign y5 = (-(^((~$signed((p12<=a4)))<=((|b2)==(+a3)))));
  assign y6 = $signed((3'd0));
  assign y7 = {4{((3'd3)>>>(^b3))}};
  assign y8 = $unsigned($unsigned($unsigned((({4{{4{a1}}}}!=(({2{a2}}!==$unsigned(a3))<<((a5)&(p10&p11))))))));
  assign y9 = (-$signed($unsigned((-$unsigned(((b1+a2)+$signed(b1)))))));
  assign y10 = (~&(~{{a0,b4},$signed(a3),(^a5)}));
  assign y11 = (((a2?p8:p16)?(5'd21):(p11?p11:p1))?(4'sd5):(-4'sd3));
  assign y12 = ((3'd0)^~(-4'sd4));
  assign y13 = (~((5'd2 * p12)>>(p8^p4)));
  assign y14 = {(b5?b3:a3),(a3?a5:p9)};
  assign y15 = (b5?a3:b1);
  assign y16 = ({(a3^~a1),{p7,p3,b4}}&&{(p3>=p7)});
  assign y17 = {{3{(-(p9>>>p8))}},{((p5?a5:a1)?(a2!==a1):(p3<=b1)),((p9?p13:p7))}};
endmodule
