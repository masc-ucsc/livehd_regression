module expression_00710(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-4'sd1);
  localparam [4:0] p1 = (~^(5'd26));
  localparam [5:0] p2 = ((4'sd1)?(3'sd3):((4'sd4)!=(2'd3)));
  localparam signed [3:0] p3 = {1{{1{(^{2{((5'd21)<<(-2'sd1))}})}}}};
  localparam signed [4:0] p4 = (5'd8);
  localparam signed [5:0] p5 = {((4'd15)===(4'd10)),((4'sd7)<=(-5'sd5))};
  localparam [3:0] p6 = ((&((|(3'd6))?(~^(5'd8)):((2'sd0)^(3'sd0))))<=(((-2'sd1)?(2'sd0):(2'sd1))?{4{(-2'sd0)}}:((4'sd1)?(-2'sd1):(-5'sd10))));
  localparam [4:0] p7 = {4{(3'd7)}};
  localparam [5:0] p8 = ({((3'd7)?(3'd0):(4'd1))}?({(4'd9),(4'd4),(-4'sd5)}+((4'd1)^(2'd3))):({(-4'sd1)}||(2'd3)));
  localparam signed [3:0] p9 = (4'd10);
  localparam signed [4:0] p10 = (((6'd2 * (3'd7))>>>(5'd10))>>(((2'sd0)==(3'sd0))==((4'd1)>>(4'sd4))));
  localparam signed [5:0] p11 = (5'd2);
  localparam [3:0] p12 = (((-3'sd1)>(4'd11))==((3'd4)>>(-5'sd7)));
  localparam [4:0] p13 = {3{(-5'sd13)}};
  localparam [5:0] p14 = {2{(-(3'd7))}};
  localparam signed [3:0] p15 = ((~|(!{((4'd2 * (5'd29))|(&(4'd12)))}))>{(~(-2'sd0)),(3'd7),(^(3'd3))});
  localparam signed [4:0] p16 = (((-4'sd0)!==(3'sd0))==={2{(4'sd6)}});
  localparam signed [5:0] p17 = ((((4'd13)?(2'd3):(2'sd0))?((4'sd1)&(3'd5)):{(4'd7),(3'd3)})>=(((4'sd7)>>>(2'sd1))?{1{(5'd8)}}:{4{(2'd0)}}));

  assign y0 = (6'd2 * (6'd2 * p14));
  assign y1 = ((3'sd1)==(a2!==b4));
  assign y2 = ($unsigned(p13)?(2'sd0):(~|p16));
  assign y3 = {{1{(5'd18)}}};
  assign y4 = (((b2|a1)<<<{4{a4}})!={(~|({b5,a3}<<(+a2)))});
  assign y5 = (a0?p11:b4);
  assign y6 = {(p0+p6),(p5),{b2,p11}};
  assign y7 = (({4{p9}}?(b5==b0):(a4<=p12))==(((a0<<<a3)-(a3!=a1))>=({2{a1}}==(a4?b5:p17))));
  assign y8 = (^(!{1{(|({3{(&a3)}}>>>{3{(!a0)}}))}}));
  assign y9 = (2'sd1);
  assign y10 = (((p2?p12:p9)<<<(p0!=p9))?(b2?p11:b2):($unsigned((a3^b2))));
  assign y11 = ((2'd0)<=(3'd1));
  assign y12 = (~&{(4'sd6),{a4,p9,p7},{p12}});
  assign y13 = ({4{a5}}&(b1^a4));
  assign y14 = (-5'sd13);
  assign y15 = ((p13?a5:p4)?$unsigned((2'd1)):$unsigned((5'sd5)));
  assign y16 = ((b1?a0:a3)?(p11?b2:p6):(a5?p0:b2));
  assign y17 = $unsigned(($unsigned(p16)));
endmodule
