module expression_00102(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({((4'd0)&&(-2'sd0)),((-5'sd6)>(4'd8))}<<<{(2'd3)});
  localparam [4:0] p1 = (&(|(!(^(~&(~|(&(^(!(-(+(+(-3'sd1)))))))))))));
  localparam [5:0] p2 = (|(~(((-(2'sd1))^~(|(5'sd8)))<<<(2'd1))));
  localparam signed [3:0] p3 = (((5'd3)+(3'sd1))<<((-2'sd0)>>(-3'sd3)));
  localparam signed [4:0] p4 = ((((5'sd7)?(-5'sd3):(2'd1))^((3'd0)||(2'd1)))&(((-2'sd1)<<<(-2'sd1))-(|(+(2'sd1)))));
  localparam signed [5:0] p5 = ((5'd11)-(-2'sd0));
  localparam [3:0] p6 = ({3{((2'sd1)?(5'd14):(5'd10))}}>>{4{((4'sd3)||(4'd8))}});
  localparam [4:0] p7 = ((~|(~&((5'd20)&&(-5'sd8))))-(+(((2'd3)<<<(5'd3))>>(+(-3'sd1)))));
  localparam [5:0] p8 = (2'd1);
  localparam signed [3:0] p9 = (-4'sd7);
  localparam signed [4:0] p10 = (~((((-5'sd13)-(5'sd10))-(6'd2 * (5'd5)))|(!{1{{3{(-5'sd12)}}}})));
  localparam signed [5:0] p11 = (-{(-(3'sd3)),{(4'd5),(4'd11)},{(-4'sd6),(-3'sd1),(2'd0)}});
  localparam [3:0] p12 = (+(~&(2'sd0)));
  localparam [4:0] p13 = ((3'd7)?{2{(-2'sd0)}}:(2'd0));
  localparam [5:0] p14 = ((4'd6)?(+(5'sd13)):(2'd0));
  localparam signed [3:0] p15 = (-((4'd2 * (5'd26))<(~^(3'd5))));
  localparam signed [4:0] p16 = (((|(-5'sd7))>((3'sd0)&(2'd0)))?((-5'sd3)?((3'd5)>(2'd3)):((2'd2)?(3'd0):(3'd4))):(((3'd3)!=(-5'sd2))?(~&(-5'sd1)):(&(5'sd10))));
  localparam signed [5:0] p17 = {1{{{2{(3'd4)}},(-5'sd4)}}};

  assign y0 = (p10?a3:p0);
  assign y1 = ((2'd1)-(5'd2 * (b1>=a2)));
  assign y2 = $signed(({{p12,a2},(b3<p13)}?{(p12?p0:p14)}:{(p4?p1:p2),(a4?b3:b4)}));
  assign y3 = (|(^p14));
  assign y4 = $signed(($signed((5'sd0))!=={(-a3),(a5>>a1)}));
  assign y5 = (2'd0);
  assign y6 = (+{4{p15}});
  assign y7 = (-(((~|p2)?(|a1):(p17?p10:b1))<(~((b5?a4:p12)|(!(p1<<p2))))));
  assign y8 = (-p7);
  assign y9 = (+{{(+p10),(-b2),{a3}},((~&p11)?(p15?p13:p9):(+p0))});
  assign y10 = (p0&&p16);
  assign y11 = ((4'd2 * (p8&a1))&&{{b0,a4,b5}});
  assign y12 = (~^((~^(~|(^{(~a3),{a1}})))&&((~^(~a5))>>(!(b2!=a1)))));
  assign y13 = ((-(p14>=p5))<<((+b2)-(~p4)));
  assign y14 = ((~^(~|(p4<=b2)))>>>((b1>>b2)===(&b0)));
  assign y15 = $signed(({(!b4),$unsigned(a0)}<<<(-$unsigned((!(~|p15))))));
  assign y16 = (({3{a3}}?(^$signed(p10)):$unsigned($signed(p15)))&(({4{p7}}?{4{p3}}:(p16))<<((p16?p3:p13)?(p3?p17:p12):(p7^~b3))));
  assign y17 = (((p4?a4:a3)>>>(p14!=p11))?((a5?p11:b2)*(b4!=b5)):(a4?p1:a3));
endmodule
