module expression_00981(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{3{(~^(4'd0))}}}};
  localparam [4:0] p1 = {{2{{(|(4'd0))}}},{3{{(3'd3),(4'sd5)}}}};
  localparam [5:0] p2 = (((3'sd0)>(-4'sd2))?((4'd5)?(4'd5):(-2'sd1)):{2{(3'd1)}});
  localparam signed [3:0] p3 = ((~^((3'd4)<<<(5'd25)))?(!((4'sd6)!==(5'd22))):((4'd15)?(4'd9):(2'd2)));
  localparam signed [4:0] p4 = (~^((((-3'sd2)|(3'd6))>>{(4'd1)})<={(-{(-2'sd0),(2'd3),(4'd0)})}));
  localparam signed [5:0] p5 = {4{(4'd13)}};
  localparam [3:0] p6 = {(!{(3'sd3)}),((5'd10)?(5'd4):(-5'sd13)),((3'd1)^~(5'd31))};
  localparam [4:0] p7 = (((((2'sd1)&&(3'sd0))+((3'd1)<(5'd19)))&((4'd2 * (5'd20))==((2'd3)!==(4'd12))))===((&((4'd11)!==(5'd2)))>(~|(~((2'd0)|(-4'sd5))))));
  localparam [5:0] p8 = (4'd2);
  localparam signed [3:0] p9 = (((2'd0)||(4'd9))>((-4'sd0)||(-5'sd12)));
  localparam signed [4:0] p10 = ((2'sd0)?((3'd4)>(-2'sd1)):((3'd0)<<<(4'd4)));
  localparam signed [5:0] p11 = (((5'sd6)?(3'd7):(5'd24))|(^((-4'sd0)>>>(-2'sd1))));
  localparam [3:0] p12 = (!(((!(-3'sd1))&&((2'sd1)+(3'd3)))&&(+(|(~^(5'sd7))))));
  localparam [4:0] p13 = (((2'd1)?(4'sd4):(-4'sd2))?((-4'sd6)?(5'sd3):(3'd1)):{(2'd0),(4'd11),(5'd21)});
  localparam [5:0] p14 = (-(((-(~|(3'd7)))/(-5'sd11))<(((4'sd1)?(5'sd5):(4'sd3))%(2'd0))));
  localparam signed [3:0] p15 = (((4'd1)<=(-4'sd3))&((5'd28)>>>(3'sd3)));
  localparam signed [4:0] p16 = {3{((4'sd1)?(2'sd0):(4'd6))}};
  localparam signed [5:0] p17 = {2{((4'sd5)?(-2'sd0):(2'd1))}};

  assign y0 = {1{{3{(p5<=a4)}}}};
  assign y1 = (((p3?p6:b5)?(p0?b2:p1):(b3|p1))||(3'd1));
  assign y2 = (~^(2'd1));
  assign y3 = ((~&(!{4{{1{p13}}}}))>$signed(($signed((p9?p8:p6))>{2{(~&a3)}})));
  assign y4 = (-(4'sd5));
  assign y5 = (((p17<=p3)+(5'd19))||$unsigned((4'd6)));
  assign y6 = (3'd1);
  assign y7 = ((^(~^b1))%a4);
  assign y8 = (~(~&$unsigned(($unsigned(({2{a3}}<<{1{$signed(b1)}}))!=={1{{3{(b2?a5:a3)}}}}))));
  assign y9 = {b1};
  assign y10 = (({b5}||(2'sd0))>=(~&(&(3'd3))));
  assign y11 = $unsigned($unsigned($signed(a3)));
  assign y12 = {{p2,p3},{p6},{p13}};
  assign y13 = (((!b4)?(p10+b0):(p7?b2:p1))||({(p10|b1)}&&{p15,p4,p12}));
  assign y14 = (4'd6);
  assign y15 = (!{((&(p15<<p16))>(p3-p14)),(+$signed($signed((-$unsigned({3{p9}}))))),$unsigned(({4{p17}}<<{p15,p16}))});
  assign y16 = {2{(5'd15)}};
  assign y17 = {b3,p4,a5};
endmodule
