module expression_00716(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(5'd8)}};
  localparam [4:0] p1 = (+((((-3'sd1)-(2'd2))>>((3'sd0)+(5'd20)))<<(~&({1{(3'd6)}}!=((-2'sd0)>>>(2'd3))))));
  localparam [5:0] p2 = ((5'd2 * {(2'd1),(5'd7),(5'd2)})===((6'd2 * (2'd2))<=((2'd2)^(5'd19))));
  localparam signed [3:0] p3 = ((~&(((4'd15)-(-4'sd4))^~(-{(-5'sd10),(2'sd0)})))+((-{(-4'sd6),(4'sd1),(3'd2)})<<((3'd0)<=(5'd30))));
  localparam signed [4:0] p4 = (~((2'd1)>({(|(5'sd10))}^(5'd19))));
  localparam signed [5:0] p5 = (!((~&((2'd3)+(-3'sd2)))+(~^(+(5'd2)))));
  localparam [3:0] p6 = (({(5'd14),(-4'sd6)}^~(3'sd0))&&(3'sd2));
  localparam [4:0] p7 = ({((4'd5)?(4'sd6):(3'd1))}=={(-4'sd2),(5'd11)});
  localparam [5:0] p8 = {4{(3'sd2)}};
  localparam signed [3:0] p9 = ((~&(3'd4))==((3'd6)<<<(-3'sd2)));
  localparam signed [4:0] p10 = ((4'd10)+(-3'sd0));
  localparam signed [5:0] p11 = ((3'd6)==={3{(-3'sd1)}});
  localparam [3:0] p12 = ((!(-(|(-(3'd3)))))>=((~&(~^(3'd1)))/(5'd8)));
  localparam [4:0] p13 = ({((-5'sd12)>(-5'sd7)),(+(3'd5)),((2'd1)?(2'd0):(3'd3))}>>>({3{(2'sd0)}}?(&(2'd3)):(~&(5'sd13))));
  localparam [5:0] p14 = {2{{{((5'sd1)?(-5'sd2):(-4'sd6)),{(-3'sd1),(5'd27)}}}}};
  localparam signed [3:0] p15 = (!(-5'sd9));
  localparam signed [4:0] p16 = (-3'sd2);
  localparam signed [5:0] p17 = {2{{1{(6'd2 * {3{(5'd18)}})}}}};

  assign y0 = ({(3'd6)}!==(6'd2 * {b2,a1,b1}));
  assign y1 = (|{((a0?a1:a5)?((2'd1)^~(2'sd0)):((a3!==b1)-(a4<<<a5)))});
  assign y2 = (-2'sd0);
  assign y3 = {p17,b3,p7};
  assign y4 = ((({1{p4}}<<<(b1<<<p5))>>({p5,a1}<(5'd2 * p0)))>={2{((p1?p3:p6)<={p17,p3,p1})}});
  assign y5 = {3{(5'sd12)}};
  assign y6 = {1{{3{a4}}}};
  assign y7 = (^({3{{3{p1}}}}?((&p7)?{3{p7}}:(~b0)):(-(p15?p14:p8))));
  assign y8 = (~^(6'd2 * (a2?b2:b1)));
  assign y9 = ((b4)?(p14/a4):(|a0));
  assign y10 = {$signed((~^($signed(a3)<=(p5!=a0)))),(+(!({p10}&&(~|p4))))};
  assign y11 = {3{p6}};
  assign y12 = {a3};
  assign y13 = (~|(~(&(5'sd4))));
  assign y14 = (~&{(2'sd0)});
  assign y15 = (({(~|p14)}==(p14&p15))^{(p6&a5),(p16||a5)});
  assign y16 = {$signed({2{a5}}),(-2'sd0),((b5^b4))};
  assign y17 = ((a2?p1:p8)>{2{p2}});
endmodule
