module expression_00064(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd0)&(-2'sd1))>(~^(3'sd1)));
  localparam [4:0] p1 = ((~|(^(-2'sd0)))/(2'd3));
  localparam [5:0] p2 = ((5'd5)<<(4'd12));
  localparam signed [3:0] p3 = ({1{({1{(3'd2)}}||((-2'sd0)==(2'sd0)))}}<<<(((5'd9)+(2'd3))?{2{(-4'sd0)}}:{2{(4'sd6)}}));
  localparam signed [4:0] p4 = ({4{(2'sd1)}}^~(-4'sd6));
  localparam signed [5:0] p5 = ((((2'd1)?(2'd2):(4'd5))?((3'd7)?(2'd3):(-3'sd3)):((2'd1)?(2'd2):(-2'sd1)))?(((5'd28)?(2'sd0):(5'd16))?((3'd7)?(2'd1):(2'd2)):((3'd2)?(2'sd0):(5'sd4))):(((-3'sd2)?(2'sd0):(2'd3))?((4'sd7)?(5'sd8):(-4'sd3)):((2'd0)?(3'd2):(2'd1))));
  localparam [3:0] p6 = (~&(~(3'sd3)));
  localparam [4:0] p7 = {(6'd2 * ((4'd7)?(3'd3):(2'd0)))};
  localparam [5:0] p8 = ((3'd3)%(3'sd0));
  localparam signed [3:0] p9 = ((2'sd1)|((3'd0)?(3'd1):(-2'sd0)));
  localparam signed [4:0] p10 = {1{({1{(-(&((-5'sd6)^~(5'd12))))}}&&{3{(-5'sd14)}})}};
  localparam signed [5:0] p11 = ((((5'd1)&(4'sd5))?((3'sd0)?(4'sd6):(5'd9)):((4'd14)<<<(-4'sd5)))>>{1{({3{(5'd2)}}==((4'sd6)>>>(3'd2)))}});
  localparam [3:0] p12 = (3'd3);
  localparam [4:0] p13 = (((2'sd1)<<<(-2'sd1))+(-2'sd1));
  localparam [5:0] p14 = (-{{((-3'sd0)?(5'sd6):(3'sd2)),(-(4'sd4)),((4'sd6)?(-3'sd1):(2'sd0))},{4{(4'd7)}},{(4'd3),(&(5'd30)),(2'sd0)}});
  localparam signed [3:0] p15 = {(4'd11),(3'd2)};
  localparam signed [4:0] p16 = ((-{(-3'sd0),(5'sd2),(-3'sd3)})?{3{((3'sd3)?(5'd16):(4'd3))}}:(-(~|{(2'd1),(2'd3)})));
  localparam signed [5:0] p17 = ({(4'd2 * ((3'd2)?(2'd1):(4'd6)))}?(((-4'sd0)<<(4'sd4))<<<{(5'd17),(4'sd2)}):{((2'd1)?(4'd4):(-3'sd0)),((2'sd1)<(3'sd0)),((-2'sd0)>>>(5'd19))});

  assign y0 = {(~((!p7)&&(p0>=p15))),(+{{b5},(+b4)})};
  assign y1 = $unsigned((3'd6));
  assign y2 = (-(~|({p15}<=(p15^~a5))));
  assign y3 = (((a3!=a5)!={b5,b4})|((b5&&p2)+(a3?p7:b4)));
  assign y4 = {(a3<a1),(b4!==b0)};
  assign y5 = (-5'sd1);
  assign y6 = (((p2&p17)?{p4,p7}:{3{p10}})?((p11>>>p4)!=(~|(p7!=p2))):((^{4{p5}})>={p7,p17,p2}));
  assign y7 = (|(-5'sd15));
  assign y8 = {2{(2'sd1)}};
  assign y9 = ({3{p6}}>=(3'd4));
  assign y10 = {2{(!$unsigned((~&(({4{b0}})))))}};
  assign y11 = {(4'd9),(p9?p2:p0)};
  assign y12 = {2{(3'sd0)}};
  assign y13 = (-4'sd4);
  assign y14 = $signed((-(~&((-$unsigned(((~|a1)!==(-b0))))|((~&(^b0))^~$unsigned((~&a3)))))));
  assign y15 = $signed({(b1!=b4),(!(p8?a3:p14))});
  assign y16 = (4'sd1);
  assign y17 = (-2'sd0);
endmodule
