module expression_00788(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd1);
  localparam [4:0] p1 = ((2'sd1)?(-3'sd2):{1{(5'd2 * (4'd12))}});
  localparam [5:0] p2 = ((((3'sd1)%(-2'sd0))?((-2'sd0)&&(-3'sd3)):(|(2'd0)))?(&((!(5'sd2))===((-3'sd3)?(-5'sd13):(2'd0)))):(~&(((3'sd1)>=(3'sd2))<<<((-3'sd0)|(3'd5)))));
  localparam signed [3:0] p3 = ({3{(2'd0)}}<={(-2'sd0)});
  localparam signed [4:0] p4 = ({((!((3'd2)!=(2'd0)))<((2'd0)!==(2'd1)))}>((&(!(-2'sd0)))>=(~((-2'sd1)==(5'd21)))));
  localparam signed [5:0] p5 = (~|{(!(4'd5)),((3'd2)?(5'd17):(-4'sd0))});
  localparam [3:0] p6 = ({(2'sd0),(2'sd1)}?{(4'd2),(5'd27),(3'sd1)}:((4'd3)!==(4'd13)));
  localparam [4:0] p7 = {1{((2'd3)&&(4'sd0))}};
  localparam [5:0] p8 = ((4'd9)?(-2'sd1):(-5'sd15));
  localparam signed [3:0] p9 = (~|(((4'sd2)?(4'd10):(-5'sd7))!=((4'd4)+(-5'sd5))));
  localparam signed [4:0] p10 = ((3'sd2)^~(5'd28));
  localparam signed [5:0] p11 = (((3'sd0)>(2'sd1))?((3'd0)^~(3'd2)):((2'sd1)<<(5'sd10)));
  localparam [3:0] p12 = ((~^{2{((4'd9)<(2'd1))}})===(!((-(|(2'sd1)))&(!((3'sd1)>>>(-4'sd0))))));
  localparam [4:0] p13 = (~&(+(~&(!(6'd2 * (-((5'd7)<<(5'd17))))))));
  localparam [5:0] p14 = (((2'sd0)?(4'd12):(4'sd5))|(^((3'sd3)<=(4'd1))));
  localparam signed [3:0] p15 = (((!(-(~^(4'd15))))<=(~|((2'sd0)>(5'd30))))-(|(~&((&((3'd3)===(3'd5)))>>>(6'd2 * (2'd3))))));
  localparam signed [4:0] p16 = (-((&{2{(-2'sd0)}})!==((2'sd1)||(5'sd0))));
  localparam signed [5:0] p17 = {{{2{(3'd7)}},{2{(5'd21)}}},{4{(-4'sd4)}},{1{{{1{(2'sd1)}}}}}};

  assign y0 = (p4?p17:p0);
  assign y1 = {4{(p9+b3)}};
  assign y2 = (((a0>>p10)*(5'd2 * p7))>=(((b4<<<a1)-$signed(a4))+((a4-b0)!==$unsigned(b5))));
  assign y3 = ({a1}||(a2<p5));
  assign y4 = ((5'sd15));
  assign y5 = (a0?a4:p8);
  assign y6 = (((+$signed(a0))>>(^(b4<<<b1)))&&((b0<b1)&&(+$unsigned(p17))));
  assign y7 = (2'sd0);
  assign y8 = $signed(((a1)?(~b2):(3'd3)));
  assign y9 = (3'd0);
  assign y10 = (2'd2);
  assign y11 = (p9^p4);
  assign y12 = ({4{b1}}-((!a1)<<<(a4!=a2)));
  assign y13 = (&(6'd2 * (p14<<<a1)));
  assign y14 = (!(4'sd3));
  assign y15 = ((p11?b3:p17)>>{(p2?p16:p13),(a0<<<p1)});
  assign y16 = {{(+p2),(~&b5)},{(b3?a0:a2),{2{p8}},{3{a1}}}};
  assign y17 = ({(((|p11)&&(p16?p16:p8))>>>(~^(!(&p11))))}|((p11?p13:p16)?(p11?p2:p15):(p14?p8:p12)));
endmodule
