module expression_00551(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(-5'sd9),(-3'sd3)};
  localparam [4:0] p1 = ((!(-((5'sd2)|(3'sd1))))==((5'd2 * (5'd4))>>((4'sd5)>=(4'd10))));
  localparam [5:0] p2 = ({4{(&(2'd1))}}&(|{4{(2'sd1)}}));
  localparam signed [3:0] p3 = (!{4{((-2'sd0)==(2'd2))}});
  localparam signed [4:0] p4 = (5'd2 * ((4'd5)!==(5'd6)));
  localparam signed [5:0] p5 = (~&((5'sd13)^(4'd12)));
  localparam [3:0] p6 = ((4'd11)==(-5'sd14));
  localparam [4:0] p7 = ((((4'sd0)?(-2'sd1):(2'd3))?(~|(3'sd0)):{2{(-2'sd1)}})+(((3'd2)?(3'd6):(-4'sd7))===(^((2'd0)>>>(3'd1)))));
  localparam [5:0] p8 = (|((4'sd3)&&(&((-5'sd1)>(5'd18)))));
  localparam signed [3:0] p9 = (-2'sd1);
  localparam signed [4:0] p10 = ((((-2'sd0)^(2'd2))?((3'sd2)?(3'd6):(5'd22)):((2'sd1)?(3'sd2):(5'd31)))?(2'sd1):((-(4'd10))?((5'd10)?(2'sd0):(2'sd0)):((5'd25)!=(-5'sd0))));
  localparam signed [5:0] p11 = {((~^(2'sd0))<<(-(5'd25))),{2{{2{(5'sd11)}}}},(((5'd21)!=(2'd0))>=((5'd14)<<<(5'sd4)))};
  localparam [3:0] p12 = (((-2'sd0)*(-5'sd2))>((4'sd5)&(5'd6)));
  localparam [4:0] p13 = {3{{4{(5'd6)}}}};
  localparam [5:0] p14 = (4'sd5);
  localparam signed [3:0] p15 = {4{(2'd0)}};
  localparam signed [4:0] p16 = ({2{(-(4'd8))}}?(4'd13):((~^(-2'sd0))>=((3'sd1)+(-5'sd10))));
  localparam signed [5:0] p17 = {2{(3'd7)}};

  assign y0 = {4{$signed(b5)}};
  assign y1 = (~|(3'd7));
  assign y2 = ((-(~^(!b0)))!=={1{{3{a4}}}});
  assign y3 = ((a1)?(5'd18):$signed(b3));
  assign y4 = (p6?b4:b3);
  assign y5 = (-(5'd27));
  assign y6 = (~|{1{{(-{(~|(2'd1))})}}});
  assign y7 = (&(&(~^$unsigned({(+(5'd6))}))));
  assign y8 = (~&(~&(~(2'd3))));
  assign y9 = ({4{(2'd2)}}>(4'sd6));
  assign y10 = ((3'd0)?(a0||p8):(a3^~p14));
  assign y11 = (($signed(((b2)>>(a3?b4:b2)))+((a0-b4)-(a1?a2:a5)))||(((b5^b2)?(b0>b2):(a5))^((b1)!==(b1?b0:b4))));
  assign y12 = (|{4{(b0?a5:b0)}});
  assign y13 = {{b2,p6,p0}};
  assign y14 = (^$signed($signed(((+p9)))));
  assign y15 = ({4{$signed($unsigned((&p13)))}});
  assign y16 = $unsigned(p0);
  assign y17 = (((6'd2 * b1)!=(-5'sd0))<={{a3},(a3&b0)});
endmodule
