module expression_00627(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{{(2'sd1),(3'd6),(4'd4)}},{(2'd2),(4'd8),(-2'sd0)},{(-2'sd0),(2'd1),(3'd0)}};
  localparam [4:0] p1 = {2{(-3'sd2)}};
  localparam [5:0] p2 = (((~|((5'd25)|(4'd13)))>>((-2'sd0)>(2'd0)))<(~^(((5'sd11)|(3'd2))>=((2'd3)&(5'd19)))));
  localparam signed [3:0] p3 = (({4{(-4'sd5)}}|(5'd2 * (3'd5)))+{4{(3'd6)}});
  localparam signed [4:0] p4 = ((((-2'sd0)>=(5'sd6))>{(5'd5),(-2'sd1),(5'd17)})===(((4'sd3)<<(-2'sd1))===((5'd27)<<(3'sd3))));
  localparam signed [5:0] p5 = ((4'd8)>>>(2'd0));
  localparam [3:0] p6 = {4{{3{(2'd3)}}}};
  localparam [4:0] p7 = ((((5'd27)!=(4'sd7))&(4'd15))?(-2'sd0):(2'd1));
  localparam [5:0] p8 = ((&({{(5'd11)}}!={(3'd7),(2'd3)}))>>>{(|(~(3'sd0))),(~|{(5'd18),(3'd4)}),(~&(!(-5'sd15)))});
  localparam signed [3:0] p9 = ((((3'sd3)?(-3'sd0):(5'sd14))&&((3'd6)+(4'd5)))?(((2'd2)?(-2'sd0):(-5'sd5))===((4'd15)?(3'd3):(-4'sd6))):((-4'sd0)?(4'sd6):(3'd3)));
  localparam signed [4:0] p10 = ((5'd24)?({(5'd3),(5'd26),(3'd2)}>{4{(2'd1)}}):(((-3'sd2)?(-4'sd0):(3'sd1))&&((3'd7)||(-2'sd0))));
  localparam signed [5:0] p11 = {2{(-5'sd2)}};
  localparam [3:0] p12 = ((((-3'sd3)===(-4'sd4))>=(4'd2 * (5'd10)))!==(((2'd1)>=(5'd20))+((-2'sd1)<(2'd1))));
  localparam [4:0] p13 = (((2'd2)>=(4'd14))<=((2'd3)/(-2'sd0)));
  localparam [5:0] p14 = {2{({1{(2'sd1)}}?{1{(4'sd2)}}:{4{(5'd12)}})}};
  localparam signed [3:0] p15 = {((((-5'sd9)|(5'sd6))>>>((5'sd2)<(-5'sd7)))>>>(((-2'sd0)!=(4'sd4))^(5'd2 * (5'd18))))};
  localparam signed [4:0] p16 = {1{(({{1{(4'd15)}}}+((5'd26)>(-5'sd2)))===((-(-(3'd4)))<=(&{4{(-4'sd3)}})))}};
  localparam signed [5:0] p17 = (~&((&(|((3'sd2)?(5'd15):(5'd15))))===(((2'sd0)?(3'd1):(-4'sd7))<<(~&(5'd28)))));

  assign y0 = {(b3<<p2),(5'd17),(-5'sd3)};
  assign y1 = (((6'd2 * (p1*a0))<<(~|(b5>>>p5)))|($unsigned((p13&&p17))<(&(p13<p2))));
  assign y2 = (^((b4/b2)+(|(^a3))));
  assign y3 = (~&(+((3'd7)^{(-4'sd7)})));
  assign y4 = $unsigned({2{(&(3'sd3))}});
  assign y5 = {({p3,p7,p11}&&(p2?p17:p15)),((&p6)?{p6,p11}:(5'd2 * p12)),(|((p6?p7:p12)==(!p12)))};
  assign y6 = (-2'sd1);
  assign y7 = (5'd15);
  assign y8 = (((b0<=p9)&(b4|p15))?((b3-a5)===(&b1)):(p9?p14:p11));
  assign y9 = {2{($signed((p13?a1:p5))?{2{a1}}:(2'd0))}};
  assign y10 = {(((p17-p1)<<<{a0,a0})+({p1}&{b1})),{{{p13,b2}},{p10,p2},(p2|p8)}};
  assign y11 = ((^p15)<<<{1{p1}});
  assign y12 = ((b1?p14:p8)?(((~&b3))):$unsigned((p4?p15:a0)));
  assign y13 = (((~&(a4?a4:a1))?(a2===b1):(~^(a0&&a3)))>>>(+(-{1{((|a2)^(6'd2 * a2))}})));
  assign y14 = (-((~^(~&$unsigned((~$signed((!$unsigned((p1?p6:p7))))))))));
  assign y15 = ((-((4'd8)>>>((4'd12)<<<(!b0))))&((+{4{a5}})!={1{({4{b5}}>>>(b0&&a5))}}));
  assign y16 = {{(p4!=a2),(p15+b0)},({((b1||a4)>(a0>>p2))}),{$unsigned(((b1||p1)^(b1)))}};
  assign y17 = {2{(~^(-{1{((p1?p14:a5)?(p8?a4:p8):(~^p7))}}))}};
endmodule
