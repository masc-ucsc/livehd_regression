module expression_00643(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd2);
  localparam [4:0] p1 = {{1{{(5'sd13),(5'd4)}}},{{4{(2'd0)}}},{{(5'sd7),(3'd3),(4'sd7)}}};
  localparam [5:0] p2 = ({((-2'sd0)?(4'd10):(-5'sd9)),((-3'sd2)!=(4'sd4))}&{((5'd9)?(-4'sd4):(4'd8)),((3'd3)&(-5'sd5))});
  localparam signed [3:0] p3 = ((~&(5'd18))?{4{(2'd1)}}:((5'sd13)?(4'd14):(-5'sd10)));
  localparam signed [4:0] p4 = ((&(+{{2{(-2'sd1)}},((2'd2)!==(3'd1)),{(3'sd0),(5'd23)}}))^(((3'sd0)?(-3'sd0):(2'd3))!=={(5'd30),(-3'sd2),(-3'sd3)}));
  localparam signed [5:0] p5 = ((~|{(2'd2),(3'd3),(5'd12)})-((~|(-2'sd0))>{(3'd4),(-2'sd0)}));
  localparam [3:0] p6 = (^(|(^((3'sd2)&&(3'sd3)))));
  localparam [4:0] p7 = {{3{{(-5'sd1),(-3'sd1),(5'd30)}}},(5'd25)};
  localparam [5:0] p8 = {{(~|((4'sd0)?(-2'sd1):(5'd24))),{(2'd0),(4'sd0),(-3'sd3)}},{(+(5'd6)),(~|(2'd0)),(!(-5'sd9))}};
  localparam signed [3:0] p9 = {((4'd1)<=(2'd2))};
  localparam signed [4:0] p10 = ((3'sd0)==((3'd7)<<(5'd9)));
  localparam signed [5:0] p11 = (((2'd2)?(2'd2):(2'sd0))?(5'd10):(2'd2));
  localparam [3:0] p12 = ((5'sd3)!==(4'd2 * ((3'd6)&(3'd5))));
  localparam [4:0] p13 = (((~&{1{(4'd2)}})>>((4'sd0)>=(3'd7)))||{(3'd5),{1{{(-2'sd0),(-2'sd0),(3'd0)}}}});
  localparam [5:0] p14 = (((-2'sd1)&((5'sd5)^~(2'sd1)))>(-5'sd11));
  localparam signed [3:0] p15 = {1{(-2'sd1)}};
  localparam signed [4:0] p16 = (5'sd15);
  localparam signed [5:0] p17 = ((((4'sd5)^~(3'd0))%(-2'sd0))>>>(((-3'sd0)<(2'sd0))^~((4'd11)+(5'd5))));

  assign y0 = (p2|p16);
  assign y1 = (4'd2 * (b0^~a0));
  assign y2 = ({1{{4{b4}}}}?{2{(-3'sd2)}}:(5'd0));
  assign y3 = (3'd6);
  assign y4 = {3{p15}};
  assign y5 = (~|(2'd0));
  assign y6 = (5'd9);
  assign y7 = (~|((a2?a1:b1)?(|{a5,b4,b0}):{(~&b1),(~a2)}));
  assign y8 = ({1{({3{p7}}==(4'd15))}}!={4{(~^p8)}});
  assign y9 = (-$signed({$signed((~((^(~&(p0)))))),({p5,a2,p11}?(p16?p16:p8):(p10))}));
  assign y10 = (~|p12);
  assign y11 = {1{{(p12|p3),{3{p12}}}}};
  assign y12 = ((+(~|{2{a3}}))?({3{a1}}<<(a0||b4)):{2{(a4==a3)}});
  assign y13 = (~((&(b5^~b3))!==(b0-b0)));
  assign y14 = {3{p16}};
  assign y15 = (-(-4'sd4));
  assign y16 = (({(2'd3),(a5<<<b2)}&(~&{b4,b5,b0}))===((4'd14)<<(+(4'sd3))));
  assign y17 = (&($unsigned({(p9>=a5)})?(+(p6?b0:b4)):((a5)>>{p12,p10,p8})));
endmodule
