module expression_00658(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{1{(4'sd3)}},{1{{(5'sd4),(4'd7),(4'd5)}}}};
  localparam [4:0] p1 = ((3'd4)!==(5'd13));
  localparam [5:0] p2 = (3'd1);
  localparam signed [3:0] p3 = (^(((3'sd3)<<<(-3'sd0))<=((2'sd0)|(5'sd6))));
  localparam signed [4:0] p4 = (~(5'd26));
  localparam signed [5:0] p5 = (^((5'sd4)>=(2'd1)));
  localparam [3:0] p6 = ((4'd13)+(-2'sd0));
  localparam [4:0] p7 = {3{((4'd13)?(5'd26):(4'sd4))}};
  localparam [5:0] p8 = ({(5'sd2),((5'd0)===(2'sd0))}?{2{(2'sd0)}}:({(5'sd6)}?(4'd12):((-4'sd2)>(3'd0))));
  localparam signed [3:0] p9 = (3'sd2);
  localparam signed [4:0] p10 = ({((-4'sd5)?(3'd1):(-3'sd0)),((3'sd2)?(4'd2):(2'sd1))}!=={({2{(4'd11)}}!==((-5'sd9)?(-4'sd7):(2'sd0)))});
  localparam signed [5:0] p11 = ((~(!((-2'sd0)>(5'd24))))==(((-2'sd1)>>>(2'sd1))<<<{2{(5'd16)}}));
  localparam [3:0] p12 = ((~|(((4'sd7)?(2'd3):(5'd5))>>((3'sd1)==(2'sd0))))>>>(~(((-4'sd0)?(2'd0):(-2'sd1))?((2'd3)?(5'd25):(3'sd0)):(~|(-5'sd15)))));
  localparam [4:0] p13 = (+{(^((!(3'sd2))?(~(4'd5)):{(2'd3),(4'd3),(5'sd2)})),({(5'd19),(-3'sd2),(2'd0)}>=((3'd2)>>>(5'sd0)))});
  localparam [5:0] p14 = ((4'sd4)>(4'sd2));
  localparam signed [3:0] p15 = (|(4'd5));
  localparam signed [4:0] p16 = (&(+(((5'd26)+(-3'sd0))>((-5'sd10)||(2'd0)))));
  localparam signed [5:0] p17 = ((((3'd1)*(2'd3))|(((-4'sd1)>>(5'd9))^~((3'sd3)||(-4'sd7))))===(3'd5));

  assign y0 = ((((b2<<b2)<<$signed(a4))<=((3'd4)||(~a0)))<<$signed($unsigned(((5'sd0)<<<(!(+$unsigned(a2)))))));
  assign y1 = (~|(&(~&{(~(~&(!({b3,p9,p12}&(!b0)))))})));
  assign y2 = (((b1?p5:b0)&&(-a0))?((b2>>>p1)%p13):((b3?b0:p13)/p10));
  assign y3 = (((4'sd5)?(p14?a4:p15):{1{p8}})>((~|p4)-{3{p16}}));
  assign y4 = (a2?a4:p11);
  assign y5 = {3{(+(3'd7))}};
  assign y6 = $unsigned((^$unsigned(p12)));
  assign y7 = (2'sd1);
  assign y8 = ((4'd5)+{(4'sd7),{a5,p11,b5}});
  assign y9 = (b0-p2);
  assign y10 = ((|$signed((a5?b3:a1)))?{1{(+$signed((b0^~b1)))}}:{(a0>>p12),(5'd31)});
  assign y11 = (4'd5);
  assign y12 = (2'd1);
  assign y13 = (((a4?a4:a3)?(b2?a1:p12):(a5))?(~^(5'd2 * (^(b1?a1:b1)))):{(a2>>>a5),((a4?p17:b3))});
  assign y14 = {2{((p16?p15:p3)>>(b2||p17))}};
  assign y15 = ((a4?b5:p11)?((p9>=p1)>=(b3?b0:p11)):(p9?p17:p2));
  assign y16 = (((~|(a2|a2))==(a0<a5))>=((b2>>b4)<<(~(-a2))));
  assign y17 = $unsigned(((^p17)^(p16)));
endmodule
