module expression_00015(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'sd6)>>(4'd6));
  localparam [4:0] p1 = ((~|((6'd2 * (3'd4))-(~&(!(-2'sd0)))))===(~|(((3'd0)>>(2'd2))|((2'd2)^~(3'd3)))));
  localparam [5:0] p2 = {1{{2{(5'sd5)}}}};
  localparam signed [3:0] p3 = ((!((5'd15)^(4'd14)))>>>(4'sd4));
  localparam signed [4:0] p4 = ((4'd3)!==((5'sd3)||((5'd22)|(5'd29))));
  localparam signed [5:0] p5 = ((^((3'd1)+(-5'sd4)))%(3'd0));
  localparam [3:0] p6 = ({1{(^({4{(-4'sd6)}}|((5'd2)&(-3'sd0))))}}<<(~(~|{2{((-5'sd11)>>>(4'sd2))}})));
  localparam [4:0] p7 = (~|(~((6'd2 * (^(3'd7)))?((5'd10)?(5'sd5):(-5'sd15)):({1{(2'd2)}}===((4'sd3)?(4'd10):(-5'sd5))))));
  localparam [5:0] p8 = {3{((-3'sd1)?(5'sd3):(-3'sd2))}};
  localparam signed [3:0] p9 = ((~(2'sd0))==((-4'sd3)^~(4'd15)));
  localparam signed [4:0] p10 = ({4{{2{(-5'sd6)}}}}>>({3{(5'd23)}}-((5'd5)!=(5'sd13))));
  localparam signed [5:0] p11 = {{(-3'sd1),(-2'sd0),(5'd18)},{{{(4'd10)}}},(&{(-3'sd0),(-5'sd13)})};
  localparam [3:0] p12 = ({{(-4'sd4),(4'd14),(5'sd4)}}>>((5'd7)?(-5'sd2):(3'd3)));
  localparam [4:0] p13 = {3{(|(~&(-{1{(5'd29)}})))}};
  localparam [5:0] p14 = (2'd1);
  localparam signed [3:0] p15 = (5'd31);
  localparam signed [4:0] p16 = (((-3'sd3)||((5'd17)?(-3'sd2):(4'sd7)))?(5'sd2):{1{({2{(-4'sd4)}}==((5'd19)?(4'sd5):(-2'sd1)))}});
  localparam signed [5:0] p17 = (+{(5'd28)});

  assign y0 = $unsigned(((6'd2 * a1)^(p2>p14)));
  assign y1 = ((((p12|p9)|{4{p10}})<=(~^((!b4)>=(p16^p1))))^~{3{(&{p11,p13,a0})}});
  assign y2 = (p15?p9:p13);
  assign y3 = ({2{(3'd2)}}^{{p2,p9,p12}});
  assign y4 = ({(p11?p9:b1),{p3}}&&((p8-p11)));
  assign y5 = {2{({(a4),{1{a1}},(3'sd3)})}};
  assign y6 = (~|p8);
  assign y7 = {((p15?b5:a0)?(a5>>a4):(b0!==b5))};
  assign y8 = (3'd4);
  assign y9 = {4{(^(!(!(|b1))))}};
  assign y10 = {{3{a3}},((2'd1)===(a4>>>b4))};
  assign y11 = (b4===b1);
  assign y12 = (4'sd2);
  assign y13 = ((p9||p12)?(p8<<p10):(p8?p5:p8));
  assign y14 = ({4{(a2?p7:b3)}}?((p2<<a4)+(a3?p10:a4)):((3'sd3)^~(b3||a1)));
  assign y15 = ((~|(&(~^(|((~|{a4,p13,b3})&&$unsigned((^(-{a2,a5})))))))));
  assign y16 = (^({1{(!(~^b3))}}?((p11<=a3)&(&a2)):{1{{(a2?p14:p9)}}}));
  assign y17 = (|((3'sd0)<((4'd2 * a1)?(b3<<<b5):{b1,a1})));
endmodule
