module expression_00991(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-(^((-2'sd1)&&(2'd3))))?(3'sd3):(~^((3'd2)?(-5'sd6):(2'd3))));
  localparam [4:0] p1 = ({4{(5'd1)}}|(5'sd2));
  localparam [5:0] p2 = (~^(~(((-2'sd0)-(5'd31))*(~((-4'sd6)*(-2'sd1))))));
  localparam signed [3:0] p3 = (3'd5);
  localparam signed [4:0] p4 = (~&(2'sd1));
  localparam signed [5:0] p5 = ((^(5'd3))<=(-(4'd10)));
  localparam [3:0] p6 = (((4'sd2)^~(5'sd5))-((-5'sd6)<=(-2'sd0)));
  localparam [4:0] p7 = ({1{{4{(4'd7)}}}}&&{2{{2{(3'sd2)}}}});
  localparam [5:0] p8 = ((((4'd10)!==(-4'sd0))<{3{(4'd8)}})>>(((2'd0)>(2'sd1))?((3'd4)?(2'd1):(-5'sd9)):((2'd0)&(-2'sd1))));
  localparam signed [3:0] p9 = ({1{(~|(-5'sd6))}}!=={4{(3'd7)}});
  localparam signed [4:0] p10 = ((((-5'sd13)+(-4'sd1))+((-2'sd0)?(3'sd1):(4'd1)))?((~(5'd3))+((-5'sd15)<<<(3'sd1))):(((4'sd4)?(5'sd15):(4'd2))?((4'd13)?(4'sd6):(2'd3)):((2'sd1)<(3'd4))));
  localparam signed [5:0] p11 = ((~&((-5'sd3)?(4'd3):(4'd8)))?((5'd10)<(4'sd5)):((3'd3)?(3'd5):(5'sd13)));
  localparam [3:0] p12 = (-(((4'd8)?(2'd2):(-2'sd0))?{1{(4'sd0)}}:(-4'sd3)));
  localparam [4:0] p13 = (5'sd12);
  localparam [5:0] p14 = {((-5'sd14)?(-5'sd14):(5'd17)),((3'sd1)?(3'd0):(3'd1)),((3'sd0)?(5'd0):(-4'sd3))};
  localparam signed [3:0] p15 = {4{(5'd25)}};
  localparam signed [4:0] p16 = (3'sd0);
  localparam signed [5:0] p17 = ({1{(5'd19)}}|((5'sd9)<<<(-3'sd3)));

  assign y0 = (-{3{({2{p16}}!=(^(!p17)))}});
  assign y1 = ((~^(p4?p10:p11))>((p17?b0:p15)<(p14?p12:p15)));
  assign y2 = {2{(((!b3)+{1{a1}})+((b1>>>a5)||(~^b1)))}};
  assign y3 = (~|(4'd9));
  assign y4 = ((~(5'd2 * (^p7)))<(-((!b5)<<<(2'd1))));
  assign y5 = ({(p14<p6),(p12|b2),(p3&p12)}<{((p7==p8)&(p1<=a3))});
  assign y6 = (5'd30);
  assign y7 = (((p6&p6)==(p5^~b4))<<((p1<=p7)>=(p13>>p12)));
  assign y8 = ((&(-2'sd1))?(~^(~^(&$unsigned(b2)))):(4'sd1));
  assign y9 = {2{(!((!(4'sd7))&(2'sd0)))}};
  assign y10 = ({1{($unsigned((b5-p15))^(a5^p16))}}<<((b4^a2)^(b3-p15)));
  assign y11 = {2{(^(p13<<p12))}};
  assign y12 = ({3{(-2'sd1)}}<<<{{2{p3}},(3'd6),{p2,p7}});
  assign y13 = ((&{4{(+b4)}})>>({4{a0}}>>>((5'sd8)||(b4===a5))));
  assign y14 = (~&(-5'sd7));
  assign y15 = {(^{(~|b2),{4{a5}},{1{a5}}}),(~^(~{p11,p3,a3})),({1{{1{{p1,a2,p3}}}}})};
  assign y16 = (~((b4>>p11)?(a2?b5:b3):(^(p5<a4))));
  assign y17 = $signed(({1{((4'd5)+(p11>p9))}}&(2'd3)));
endmodule
