module expression_00876(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd1)^(4'sd5))<<((-3'sd0)?(3'd0):(5'd17)));
  localparam [4:0] p1 = (|((~(-(2'sd0)))?(!(4'd10)):(~|((3'd3)?(2'd1):(5'd12)))));
  localparam [5:0] p2 = ((2'd1)<(4'sd3));
  localparam signed [3:0] p3 = (((4'd12)==(5'd10))<(&(^(3'sd2))));
  localparam signed [4:0] p4 = ((((4'd11)>(3'd3))+(^(2'sd1)))!=={(+(3'sd0)),(~^(4'sd3))});
  localparam signed [5:0] p5 = {3{(((4'd1)<<(-4'sd0))?((3'd1)&&(5'd10)):((-4'sd2)-(5'sd6)))}};
  localparam [3:0] p6 = (2'd2);
  localparam [4:0] p7 = (-(4'd2 * (4'd8)));
  localparam [5:0] p8 = ((((5'sd8)!=(5'sd4))==={(3'd5),(2'd0),(4'd14)})+({(5'sd12),(3'd7)}!=(6'd2 * (3'd5))));
  localparam signed [3:0] p9 = (((3'd1)?(-5'sd11):(-3'sd3))?((3'd7)?(2'd3):(5'd22)):(~^((-5'sd14)?(2'sd1):(-3'sd3))));
  localparam signed [4:0] p10 = ((((3'd6)<<<(5'sd15))|((4'd12)||(3'sd2)))-(((3'd0)<<<(2'sd0))!==((4'd14)===(-3'sd2))));
  localparam signed [5:0] p11 = (!(((5'd15)?(3'd4):(4'd6))?(-((-4'sd0)?(3'd0):(5'd1))):(^((5'sd9)?(3'd1):(3'sd0)))));
  localparam [3:0] p12 = (-5'sd7);
  localparam [4:0] p13 = (-(((-5'sd6)!==(5'd12))!==((&(-3'sd0))===(5'sd9))));
  localparam [5:0] p14 = (|(({(4'd15),(-3'sd2),(2'd1)}?(^(5'sd4)):(+(2'd3)))?(~^(((2'd2)<<(2'sd1))>(~(-3'sd2)))):(~^((-(4'sd2))+(-(5'd3))))));
  localparam signed [3:0] p15 = {(+{{(5'sd11),(3'd4)},(|(~^(4'sd4))),(&(^(5'd6)))})};
  localparam signed [4:0] p16 = (((5'sd5)?(2'd1):(2'd1))>=((-4'sd7)?(4'd7):(4'sd2)));
  localparam signed [5:0] p17 = (4'd2 * (^{(5'd4),(4'd6),(3'd7)}));

  assign y0 = {{4{p16}},(p16<<p6),(&(p13&a2))};
  assign y1 = (!(!((+(+((&p16)?(~&p16):(^b5))))>((+(p10^~p7))?(p12%p7):(p3?p14:p4)))));
  assign y2 = (-4'sd0);
  assign y3 = $unsigned($signed($unsigned({{{$signed(p4),$unsigned(a2)},($unsigned($signed(p12)))}})));
  assign y4 = {{(-2'sd1),{1{{p15,p0}}},(-2'sd1)}};
  assign y5 = {2{((~^b5)!=(a1?a1:a2))}};
  assign y6 = (5'd19);
  assign y7 = ((+(~((~|(~|p0))?(^(p0?p14:p13)):(p1?p4:p3)))));
  assign y8 = (b0<<<a0);
  assign y9 = (^((&p3)=={3{a3}}));
  assign y10 = {(+(~|(5'd6))),(+{(^b1),{p6,b5,p10}})};
  assign y11 = (a1==p15);
  assign y12 = (2'sd1);
  assign y13 = (p2?a3:p14);
  assign y14 = ((((b5?b2:a0)==={1{{4{b4}}}})!=={4{(a3?a3:b2)}}));
  assign y15 = {3{{1{{4{p3}}}}}};
  assign y16 = (^(-a1));
  assign y17 = (((~|p11)?(a0*p4):(p9?p16:p3))?(~^$unsigned(((p11?p1:p5)))):$unsigned($unsigned((p1^b4))));
endmodule
