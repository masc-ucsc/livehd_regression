module expression_00284(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-5'sd8)?(5'd14):(4'd3))%(-4'sd6));
  localparam [4:0] p1 = (!(&(~(+{((3'd7)^~(5'd25)),{(5'd14),(2'd3),(5'sd9)},(&(2'd1))}))));
  localparam [5:0] p2 = ({3{{4{(-5'sd2)}}}}>>(({4{(-4'sd1)}}&(|(4'd5)))<<<((~|(5'd26))<<<{2{(-5'sd1)}})));
  localparam signed [3:0] p3 = {{(~|((2'sd1)?(2'd1):(4'd5)))},{2{((3'sd2)===(2'd3))}}};
  localparam signed [4:0] p4 = {(&(~{4{(4'sd5)}})),(!(^{{(5'd6)},(!(3'd2))}))};
  localparam signed [5:0] p5 = (4'd2 * ((5'd10)?(2'd0):(4'd14)));
  localparam [3:0] p6 = (((3'd2)!=(3'd2))?{(-5'sd12),(5'sd2),(3'sd1)}:((-5'sd14)<(-2'sd0)));
  localparam [4:0] p7 = (((5'd2)<(5'd16))&((2'sd0)%(5'sd11)));
  localparam [5:0] p8 = ({3{{(4'sd1),(-5'sd5),(2'd3)}}}>>>{{((2'd1)|(3'sd0))}});
  localparam signed [3:0] p9 = (((2'sd0)-(5'd18))<<<((-2'sd0)&&(4'sd5)));
  localparam signed [4:0] p10 = ((5'sd13)?(4'd11):(-4'sd3));
  localparam signed [5:0] p11 = (-(5'd9));
  localparam [3:0] p12 = ((4'd2 * (2'd2))===((4'sd2)&&(-4'sd7)));
  localparam [4:0] p13 = ((-3'sd1)?(4'd11):((-4'sd6)+{4{(2'sd1)}}));
  localparam [5:0] p14 = ((3'd1)===((2'd3)-(-5'sd14)));
  localparam signed [3:0] p15 = (-2'sd1);
  localparam signed [4:0] p16 = {3{((3'd7)<<(3'd0))}};
  localparam signed [5:0] p17 = {2{(5'd13)}};

  assign y0 = (~^p2);
  assign y1 = {p11};
  assign y2 = ((~^(b4))>>{p2,p10,p17});
  assign y3 = {2{{2{(5'sd11)}}}};
  assign y4 = ((&(p9>=b0))%b5);
  assign y5 = (-({3{(^a3)}}<=(!(4'd12))));
  assign y6 = (~|(3'd6));
  assign y7 = ((p4<<p12)&&(4'd2 * p13));
  assign y8 = ((&{4{(p7?p9:p11)}})?((p8)?{1{p15}}:$signed(p14)):$unsigned($signed(((p11?p15:p0)?{1{p17}}:(p17?p14:p0)))));
  assign y9 = ((p13?p15:b3)!=(b4?a0:a4));
  assign y10 = (!(~(((p10+p0)>=(p3<<<p14))<((b4>>b1)<=(b4%b5)))));
  assign y11 = (-(^((p13?p2:p5)?{p3,p10,p8}:$unsigned(p13))));
  assign y12 = (~|((~|((|b1)-(3'd5)))<=(+(~|{(!p6)}))));
  assign y13 = {{3{{1{{{1{(+{4{p7}})}}}}}}}};
  assign y14 = {2{{b3,b3}}};
  assign y15 = (!p0);
  assign y16 = (~|(4'd12));
  assign y17 = {$signed({(a2!==a3),(p17)}),(((a1^a2)===(b5|a2))),{{p14,b4,p16}}};
endmodule
