module expression_00588(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|((5'd0)<(-(-5'sd12))));
  localparam [4:0] p1 = ((+(5'sd3))<<<((!(-4'sd5))<<<((4'd11)-(3'sd2))));
  localparam [5:0] p2 = (~((-3'sd3)&(4'sd3)));
  localparam signed [3:0] p3 = (~&(~(!(~^(((-4'sd4)?(3'd6):(3'd6))?((-3'sd3)?(3'd3):(4'sd6)):(+((-4'sd5)?(4'sd1):(2'sd0))))))));
  localparam signed [4:0] p4 = {((4'sd0)?(4'd9):(-3'sd2)),{4{(5'd10)}},{(3'd1),(5'sd10),(3'sd1)}};
  localparam signed [5:0] p5 = ((2'sd1)?(2'd1):(3'sd2));
  localparam [3:0] p6 = (|(^(5'd2 * (2'd3))));
  localparam [4:0] p7 = (3'd0);
  localparam [5:0] p8 = (^((~&((5'sd5)&&(5'sd15)))===(((3'sd0)===(3'sd3))&((-2'sd0)!==(4'd14)))));
  localparam signed [3:0] p9 = (((+(&(3'sd3)))!=(+((4'd9)&&(4'd5))))>>(^((-(5'sd15))||((3'd4)==(2'd3)))));
  localparam signed [4:0] p10 = (~((2'd1)?(5'sd2):(5'd6)));
  localparam signed [5:0] p11 = (^(2'd2));
  localparam [3:0] p12 = {2{({4{(-2'sd1)}}||((-3'sd3)?(5'd5):(5'sd1)))}};
  localparam [4:0] p13 = {4{(4'd11)}};
  localparam [5:0] p14 = {3{({4{(4'd9)}}?(5'd2 * (5'd26)):(~|(3'd0)))}};
  localparam signed [3:0] p15 = {{4{{(5'sd0),(4'd7)}}}};
  localparam signed [4:0] p16 = (^((~|(6'd2 * (2'd0)))?{(-5'sd2),(5'd27)}:((4'sd3)!==(-2'sd0))));
  localparam signed [5:0] p17 = {((-(-5'sd5))?((4'sd4)?(-5'sd12):(5'd8)):((5'd18)?(5'd6):(4'sd5))),{{(2'd2),(-5'sd0)},((-2'sd1)?(-4'sd7):(2'd3))},(((5'sd10)<(4'd0))^~{(5'd19),(-2'sd1),(4'd3)})};

  assign y0 = {3{(p5?p10:p3)}};
  assign y1 = ((-5'sd9));
  assign y2 = $unsigned((((p4+p9)?(p3<=p4):(a3^p13))+({p11,a3,p1}?(3'd0):(p15&p12))));
  assign y3 = {3{{4{a0}}}};
  assign y4 = (5'd20);
  assign y5 = (-(~^(-(((~|p2)&(p15>>p9))?((b4*p2)<=(p8/p10)):((+p10)||(+p1))))));
  assign y6 = ((b4?a0:p13)^(~^{a2}));
  assign y7 = (|{2{{2{$unsigned((~(2'd3)))}}}});
  assign y8 = (((~^(6'd2 * p7))<<<((p13>=b0)-(!b3)))&((+(|b1))*(~|(p17&b1))));
  assign y9 = (({(a3==p7),(5'd2 * p0)}!={(p0<<p14)})&&{$unsigned(((p7-b3)||$signed((6'd2 * p12))))});
  assign y10 = (&(4'd2 * b1));
  assign y11 = {((b4|b3)!=(a4!==a5)),{((b5<=b5)==(a5!==a5))},({b2,a1,a3}?(a1&b4):(b4<<<b0))};
  assign y12 = ((2'd0)<=({b0,p8}?$signed(p2):{4{p8}}));
  assign y13 = {3{p2}};
  assign y14 = (~|(~&$unsigned({$signed((|$signed((!{$signed({a0,a0}),$unsigned({a3,a0,b3})}))))})));
  assign y15 = (4'd7);
  assign y16 = (((4'd2 * (b0>>a2))+(^(p1>>>p14)))>>>(~|({{p10},(~|p7)}!=({p8,p17,p10}>={p17}))));
  assign y17 = ({1{a0}}+(5'd2 * b0));
endmodule
