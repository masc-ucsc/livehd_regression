module expression_00857(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{((-2'sd0)-(3'd2))}}+({1{(6'd2 * (4'd15))}}-{2{(-2'sd0)}}));
  localparam [4:0] p1 = (2'sd1);
  localparam [5:0] p2 = {4{(4'sd4)}};
  localparam signed [3:0] p3 = ((3'd2)?(2'd0):(4'd13));
  localparam signed [4:0] p4 = {4{(&(-5'sd10))}};
  localparam signed [5:0] p5 = (~(5'd5));
  localparam [3:0] p6 = (+(-(&(5'd0))));
  localparam [4:0] p7 = (2'd3);
  localparam [5:0] p8 = (2'd3);
  localparam signed [3:0] p9 = ({((~&(3'sd3))>=((4'sd1)>(2'd3)))}>>(((-2'sd0)===(4'd6))<<{(3'd3)}));
  localparam signed [4:0] p10 = (3'd5);
  localparam signed [5:0] p11 = ((((-3'sd1)==(5'd24))>=((2'd0)%(-5'sd1)))!=(((-4'sd3)>=(2'sd0))||((2'sd1)==(3'sd2))));
  localparam [3:0] p12 = (^{(&{((4'sd1)?(2'sd1):(2'sd1)),((3'd3)>>>(3'sd2))})});
  localparam [4:0] p13 = (+(~|(|(~^(^(&(~(~^(~|(-(^(~|(5'd14)))))))))))));
  localparam [5:0] p14 = (((2'd2)?(4'd5):(4'd5))/(4'd8));
  localparam signed [3:0] p15 = {(2'd3),(3'd6)};
  localparam signed [4:0] p16 = {2{(&(-5'sd7))}};
  localparam signed [5:0] p17 = ((5'sd0)!==(2'd3));

  assign y0 = ((+(~|(((&a0)||(p1<<<a0))+((-p10)&(b2<<b1)))))<(((b1-b1)>=(p0>>b5))||(~((~b5)^(&a4)))));
  assign y1 = $signed({((2'd2)?(4'd12):(!a4)),((p17|a2)?(5'd14):(p1>=p9)),((p12>>>p3)<=$signed(b4))});
  assign y2 = {a3};
  assign y3 = ($unsigned(($signed($unsigned(p8))<(p9%p6)))&&((+(~&p10))>>>(p5||a2)));
  assign y4 = ($signed(({b0,b0}?{b5,a0}:$unsigned(b5)))!=={2{{1{{a3}}}}});
  assign y5 = {3{({4{p6}}|(b2>=p16))}};
  assign y6 = $unsigned($signed(($unsigned((p5^~b4))>>>$signed((p10^~p4)))));
  assign y7 = {3{(3'd7)}};
  assign y8 = (2'd3);
  assign y9 = ((|a1)?(-p15):(a5?a5:b4));
  assign y10 = ((a4>>a1)%a2);
  assign y11 = {4{(b4!==b2)}};
  assign y12 = (((-4'sd1)+(4'd2 * p13))+(5'd29));
  assign y13 = (|((4'd2 * (a0-b0))!==((b0>>>a0)<<(~&a1))));
  assign y14 = {$signed(p0)};
  assign y15 = {p9};
  assign y16 = (p4%b4);
  assign y17 = $signed((~(-3'sd3)));
endmodule
