module expression_00514(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(5'sd14));
  localparam [4:0] p1 = ((((5'd6)<<(3'sd2))<<<((3'sd3)%(3'sd2)))>=(((-4'sd1)<=(4'd8))===((5'd22)<=(4'sd5))));
  localparam [5:0] p2 = ((((5'd21)>(4'd4))!=={4{(5'd16)}})<=(-5'sd1));
  localparam signed [3:0] p3 = ((((5'd29)>>>(4'sd6))^((5'd16)<(5'sd10)))<<<(-3'sd2));
  localparam signed [4:0] p4 = (((-5'sd6)^~(2'sd0))?((3'd7)<<(-2'sd1)):((4'd3)?(-5'sd13):(-4'sd2)));
  localparam signed [5:0] p5 = ({((5'd27)?(-2'sd1):(4'd6))}?((4'd10)?(2'd0):(5'd7)):(2'd3));
  localparam [3:0] p6 = {(4'd2),(5'd14)};
  localparam [4:0] p7 = (|{4{{4{(3'sd1)}}}});
  localparam [5:0] p8 = (~({(2'sd0),(3'sd2)}>=(~|(-2'sd1))));
  localparam signed [3:0] p9 = {2{{3{((-2'sd0)==(4'sd7))}}}};
  localparam signed [4:0] p10 = ((5'sd12)&&(5'd3));
  localparam signed [5:0] p11 = {{(-2'sd0),(4'sd5)}};
  localparam [3:0] p12 = {3{{3{(4'd12)}}}};
  localparam [4:0] p13 = ((~^((2'sd1)!==(-5'sd15)))*((3'd2)?(4'd13):(5'd6)));
  localparam [5:0] p14 = ({3{((5'sd2)^(-5'sd0))}}<(((5'd29)|(-2'sd1))?((2'd0)?(-2'sd1):(4'sd0)):(6'd2 * (3'd0))));
  localparam signed [3:0] p15 = (((-4'sd7)?(-4'sd1):(4'sd0))>={2{(-3'sd2)}});
  localparam signed [4:0] p16 = (-3'sd2);
  localparam signed [5:0] p17 = (5'd2 * (5'd13));

  assign y0 = ({4{b1}}&(({4{b2}})));
  assign y1 = (|$unsigned(((|$unsigned(((+(-(~|$unsigned($unsigned(p11)))))||((~^$signed(b5))^~(b4===b2))))))));
  assign y2 = (!(~^(5'd5)));
  assign y3 = $signed($signed(p16));
  assign y4 = ((b1<=p16)^{p15,p16});
  assign y5 = ((((b4||b1)&&(a2))===($signed((b2>b4))))||$unsigned(($unsigned((p5^~b2))<<<$signed((b4<<a2)))));
  assign y6 = {(((|p3)?(b5!=p16):{p2,b0,b2})||{(p17?p16:b4),{2{a2}},(p13?b4:p15)}),(3'd5)};
  assign y7 = (&(~&{3{(2'd3)}}));
  assign y8 = (((!p8)?(a5!==a4):(~|p7))?((~^(~|p14))==(~(|p14))):$signed((&((~p13)|(p12>>>p8)))));
  assign y9 = ((((b4===b0)-(b3^p16))>>((p7==b1)!=(p6+a5)))==((a5&b0)?(b4===b0):(-(b3?a4:b3))));
  assign y10 = (((a2^~p16)==(|p16))<=(~(p8>=b3)));
  assign y11 = $signed({3{$unsigned($signed(p12))}});
  assign y12 = {2{b5}};
  assign y13 = ((~|(b1?p0:a4))==(-2'sd0));
  assign y14 = (6'd2 * $unsigned((p10?p15:p9)));
  assign y15 = (5'd24);
  assign y16 = {4{p9}};
  assign y17 = (+(-4'sd3));
endmodule
