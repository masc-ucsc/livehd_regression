module expression_00399(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd1)+(5'd29))+((5'd5)?(3'sd0):(3'sd1)));
  localparam [4:0] p1 = ({((2'd0)?(5'd14):(5'd18)),{(2'd1),(2'd3),(2'd0)},((5'sd15)?(4'd0):(5'sd13))}?{{(-4'sd0)},{(5'd11),(-4'sd3)},((5'd1)?(4'd5):(5'd27))}:({(2'd3),(5'd9)}?{(-2'sd1),(3'd1),(2'sd1)}:{(3'd0)}));
  localparam [5:0] p2 = (!((&{(5'sd14)})!=(^(&(4'd14)))));
  localparam signed [3:0] p3 = ({((4'd4)?(4'd8):(2'sd1)),((4'sd4)?(5'd23):(5'sd2))}?{((3'd6)?(3'd7):(5'd31)),{(2'sd1),(2'd2)},{(4'sd0)}}:{((2'd2)?(2'd3):(3'd7)),{(3'sd3),(2'sd0)},{(-2'sd0),(3'd5)}});
  localparam signed [4:0] p4 = ((~^(2'sd1))?{(-5'sd0),(2'sd0)}:{(3'sd1),(-2'sd0)});
  localparam signed [5:0] p5 = ((^((~|(-3'sd1))?(+(2'd1)):((2'd2)>(-2'sd1))))===((~^(2'd0))?(&(3'd7)):((3'd2)?(5'd16):(-4'sd3))));
  localparam [3:0] p6 = ((5'sd11)||(2'sd0));
  localparam [4:0] p7 = (((5'sd2)==(2'd0))<<<(-5'sd4));
  localparam [5:0] p8 = ((((5'd15)<(2'sd0))===((3'd3)<=(2'sd1)))+(((-5'sd0)&&(2'd1))!=={(5'd27)}));
  localparam signed [3:0] p9 = ((5'sd8)>(4'd10));
  localparam signed [4:0] p10 = {1{({2{(-3'sd3)}}?((3'sd1)<=(5'd0)):{1{(5'd2)}})}};
  localparam signed [5:0] p11 = (!(-((3'd3)<<(2'd3))));
  localparam [3:0] p12 = (~^((6'd2 * (3'd2))||(^{(2'd1)})));
  localparam [4:0] p13 = ((((-3'sd1)-(2'd3))===((4'sd4)>>(5'd19)))>=(((3'd7)<<<(3'sd0))*((3'd3)==(-5'sd14))));
  localparam [5:0] p14 = {(((3'd5)?(3'd2):(2'd0))?(~{2{(4'sd3)}}):((2'd3)?(2'd0):(4'd14))),(&{1{{4{{2{(2'sd0)}}}}}})};
  localparam signed [3:0] p15 = (~|(~|((&((2'sd1)===(3'sd2)))^{(-3'sd1),(3'sd3),(-5'sd8)})));
  localparam signed [4:0] p16 = ({{(2'd1),(4'd13),(3'sd0)}}<({(4'd14),(4'd3),(2'd2)}<((3'd5)+(-3'sd2))));
  localparam signed [5:0] p17 = (^(({3{(3'd4)}}^(!(-2'sd0)))>>{2{(~^(5'd20))}}));

  assign y0 = {({p6,p16}?{3{p16}}:(b1?p10:p14)),({a2,p2,p17}?(4'd12):(5'd25)),(~{4{p0}})};
  assign y1 = {4{{1{{3{b5}}}}}};
  assign y2 = ($unsigned((((p14<<<p1)^(b5-p0))))||(((p7^~p5))&&((p1?p17:p3)&(p1?p12:p17))));
  assign y3 = (~&(!(|(2'sd0))));
  assign y4 = (!(((~(!b2))||(b3==a2))&&{(3'd0)}));
  assign y5 = {1{($signed($unsigned($unsigned({3{(b4<<a4)}})))>>>{3{$unsigned($signed(p16))}})}};
  assign y6 = (((b2?b5:a2)==(b5?a4:a2))?((a3?a0:b0)?(a2*a2):(b4?b1:b3)):((b1==b3)?(b0+b5):(a4?b1:b5)));
  assign y7 = (^(~&(-(p16||a0))));
  assign y8 = {({p2,p12,b5}>>>{p1,a2,a3}),((!b4)<={p0,p11})};
  assign y9 = (~^(2'd2));
  assign y10 = $unsigned(($signed((~^(!p9)))?((~&a4)!==(!b5)):$unsigned({1{(~^a0)}})));
  assign y11 = $unsigned((p14?a3:p14));
  assign y12 = {2{(5'd2 * (p6&&p12))}};
  assign y13 = ({2{{1{(b1&&a3)}}}}+({4{p10}}>{3{b0}}));
  assign y14 = (((((b5)^(4'sd7))+{2{(a0)}}))-((a1&&a3)?(b4-b4):(-4'sd0)));
  assign y15 = ({3{{b2,b5}}}==={4{(b1<=b3)}});
  assign y16 = (-5'sd12);
  assign y17 = {3{{(-p3),{b0,p8}}}};
endmodule
