module expression_00214(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (6'd2 * (5'd2));
  localparam [4:0] p1 = {2{{3{(3'sd2)}}}};
  localparam [5:0] p2 = (3'd3);
  localparam signed [3:0] p3 = {({(2'sd0)}>>{(-3'sd1),(5'd27)}),(^(+{(3'd0),(4'sd7),(4'sd6)}))};
  localparam signed [4:0] p4 = (!(|{(+{((4'sd4)==(-2'sd0)),((5'd21)^~(2'd2))}),(((5'sd3)>(4'sd2))|(&(-5'sd2)))}));
  localparam signed [5:0] p5 = (!(({4{(3'd5)}}||{3{(4'd13)}})^(^{1{(5'd2 * (5'd15))}})));
  localparam [3:0] p6 = ((3'd0)==(5'sd9));
  localparam [4:0] p7 = (&{((-2'sd1)?(4'd7):(4'd13))});
  localparam [5:0] p8 = {3{{4{(2'd2)}}}};
  localparam signed [3:0] p9 = ({1{(((4'd8)||(2'd1))>>>((4'd12)!=(-3'sd1)))}}>(((2'd1)!=(2'sd1))+{4{(4'd5)}}));
  localparam signed [4:0] p10 = {4{(+{(2'sd1)})}};
  localparam signed [5:0] p11 = {(4'sd0),(5'd21),(-3'sd2)};
  localparam [3:0] p12 = {3{(+{2{{1{(-3'sd0)}}}})}};
  localparam [4:0] p13 = (((4'd6)&(-5'sd2))||((-2'sd1)<=(2'd3)));
  localparam [5:0] p14 = (-(&(3'sd1)));
  localparam signed [3:0] p15 = (((4'd8)!=(3'd0))-((3'd5)===(2'sd0)));
  localparam signed [4:0] p16 = (~{4{(4'd13)}});
  localparam signed [5:0] p17 = ({((5'd4)||(-4'sd6)),((2'd3)>(-5'sd15))}==((&{1{(5'd14)}})=={(3'sd2),(4'd11)}));

  assign y0 = $unsigned({2{$signed({1{{2{{p8,p16}}}}})}});
  assign y1 = (((a0||a4)<<(b3-a5))===((b2&a3)-(b0>a2)));
  assign y2 = ((((p11>>b4)<=(p8%a2))==((a1<=a0)<(a3<b5)))<=(((a1<=a5)<(a3%a4))^~((a3===a4)%b4)));
  assign y3 = ((a4?a0:b4)?(|(-(p14?p0:p6))):(3'd7));
  assign y4 = ((2'd3)<<((6'd2 * p12)>={b5}));
  assign y5 = (($signed({a1,a1})^~(-5'sd5))>(~&({a4,b0,b1}?(p8-b1):(a2||a1))));
  assign y6 = ({(!{b2,b3,b4}),(b1?a5:b0)}|({(4'd2 * b0)}!=(2'sd0)));
  assign y7 = (-($signed((((~^a0)<=(|a3))&{a5,b2,b5}))^~(((b4)>>>(a3&b3))=={(b1>>a3),{3{b5}},(p5<a3)})));
  assign y8 = $signed(((b3?a3:p14)?$unsigned(b1):(b2^a5)));
  assign y9 = $unsigned((-4'sd6));
  assign y10 = ((p17<<<p7)?{1{(p7>>p16)}}:(p12?p15:p17));
  assign y11 = {(((a2?a3:a0)&((a1<<a3)>>>(p10>=b0)))^~({$unsigned((b3!=b3))}>=((a2===b1)-(2'd0))))};
  assign y12 = {1{$signed({({4{{p8,a1}}}),(({2{{p4}}}||$unsigned((p9>=p16))))})}};
  assign y13 = (-(~&(~|((5'd13)?(-3'sd0):(5'd5)))));
  assign y14 = {((4'd2 * b2)!==(a5<<<a1)),({p9}<<(p0!=a2))};
  assign y15 = {b1,b0};
  assign y16 = {(p12?p5:p4),(p15?a3:p0),(b4?a5:p12)};
  assign y17 = (!(2'd2));
endmodule
