module expression_00818(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+{((-5'sd0)==(-2'sd1))})?((!(5'd9))?(~^(3'd6)):((4'sd5)-(3'd4))):((~|(3'sd2))?((-5'sd6)==(-3'sd1)):((3'd2)-(5'd14))));
  localparam [4:0] p1 = (((3'sd2)?{(4'd10)}:{4{(2'd0)}})==(((-4'sd6)>(3'd1))?((2'd0)?(3'd3):(5'sd5)):((-2'sd0)>(-3'sd3))));
  localparam [5:0] p2 = (2'd3);
  localparam signed [3:0] p3 = (((4'd10)||(-2'sd0))?(~|(!(2'd2))):((5'd26)?(5'd21):(3'sd3)));
  localparam signed [4:0] p4 = {(((2'd1)+{(-4'sd2)})?(3'd6):((2'd2)!=((-3'sd3)?(4'sd5):(-5'sd9))))};
  localparam signed [5:0] p5 = {(((~^{(-4'sd5)})<=(~|(~&(2'd2))))<<{1{(&{2{(!(2'd3))}})}})};
  localparam [3:0] p6 = ((!(4'd2))?(5'd2 * (3'd3)):((3'sd3)?(4'd11):(5'sd3)));
  localparam [4:0] p7 = {{{(3'd7)},{(4'sd5),(5'd2)}},((4'd7)?(5'sd10):((5'd0)?(4'sd5):(2'd3))),({(3'sd1)}?{(-4'sd7)}:{(2'd2),(2'd2),(5'd14)})};
  localparam [5:0] p8 = {2{({(3'd3)}<=((5'd24)>=(4'd7)))}};
  localparam signed [3:0] p9 = (3'd7);
  localparam signed [4:0] p10 = (((-3'sd2)<=(3'sd3))^(+(5'sd2)));
  localparam signed [5:0] p11 = {(5'd14),(5'd2),{({(-4'sd5),(5'd28),(5'd26)}<(~(-4'sd6)))}};
  localparam [3:0] p12 = {3{{(2'sd0),(5'sd0)}}};
  localparam [4:0] p13 = {(((4'd9)?(5'd8):(-4'sd4))?{(4'd9),(4'sd7),(5'd3)}:((4'sd5)?(5'sd12):(-4'sd2))),(5'd2 * (^{(3'd7),(4'd9)}))};
  localparam [5:0] p14 = {(-{{(~^{(-2'sd1),(5'd14),(-2'sd1)})},((~^(5'sd9))>>>{(2'sd1),(3'd4),(-2'sd0)}),({(3'd0)}==={(3'd3)})})};
  localparam signed [3:0] p15 = {4{((2'd2)+((2'sd1)!=(5'd20)))}};
  localparam signed [4:0] p16 = {4{(2'd2)}};
  localparam signed [5:0] p17 = {2{({4{(3'd0)}}|(((-3'sd3)&&(-5'sd1))+((-5'sd11)>(4'sd6))))}};

  assign y0 = ((((a0?a0:b2)>>(a5?b3:b4))+(~(b3>>a3)))==={4{(~|b5)}});
  assign y1 = {1{{(+({4{a0}}>>>(3'sd0))),{((~&p2)<$unsigned(b4))},(~^(5'd11))}}};
  assign y2 = (~|(-2'sd1));
  assign y3 = (4'd7);
  assign y4 = {((p2>>p17)>>>(p16-p1)),{(p9<p16),(5'd28),(p8&p16)},$signed(({p6,p9}))};
  assign y5 = {(5'd2 * (p0^~p6)),(({a4,a4}!={p17})>>>{(p9&&a4)})};
  assign y6 = {3{{p15,a3}}};
  assign y7 = (~^((((|b5)^~(~^a5))<=(!{{b4,b1,p17}}))>>((-((~&a3)>>(a0==a5)))<<<(!(~&(b1>=p13))))));
  assign y8 = {3{(~&$unsigned({p2,p14,p16}))}};
  assign y9 = ((~|(~|((-(a1^a4))||{3{a2}})))===(+{1{((~^(2'sd0))|{1{(b1-a0)}})}}));
  assign y10 = {{2{p12}}};
  assign y11 = (-(-b2));
  assign y12 = (((b3?b5:b4)?(-3'sd2):{b5,a3,b2})===((a5?b4:b4)?(5'd2 * b1):{{b0}}));
  assign y13 = (+($unsigned(b2)));
  assign y14 = (({{p1}}>(p2>>a3))==({(+a1)}>(b3!==b3)));
  assign y15 = (({1{((a4!==b0)^~(a1?b2:b0))}})?((a4<<<b3)?(6'd2 * b2):(a0===a1)):$unsigned({4{p16}}));
  assign y16 = ((p3?b5:p14)?(a3?b2:p3):(p10?p3:b0));
  assign y17 = (({a2,a4}===(!(a3?a4:a2)))&&(3'sd2));
endmodule
