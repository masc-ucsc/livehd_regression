module expression_00615(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(-(3'sd2))}};
  localparam [4:0] p1 = ((~|(-2'sd1))?((4'sd4)<<(3'd4)):((-3'sd0)^(5'sd1)));
  localparam [5:0] p2 = ((5'd21)?(-3'sd3):(3'd0));
  localparam signed [3:0] p3 = ({((-2'sd0)>>>(3'sd3)),{(2'd3)},(^(4'd13))}+(((-4'sd0)!=(-4'sd7))>>>{(4'sd3)}));
  localparam signed [4:0] p4 = (((3'd3)<=(-4'sd2))&((5'd29)*(4'd6)));
  localparam signed [5:0] p5 = (^((((3'd3)*(-2'sd0))?(~|(5'd29)):(~&(5'sd1)))!==(((2'd2)?(-2'sd0):(3'd3))<=(~|(-(2'sd1))))));
  localparam [3:0] p6 = {4{((4'd1)>>(5'sd9))}};
  localparam [4:0] p7 = ((+(~(-2'sd1)))>>>((3'sd0)>(4'd6)));
  localparam [5:0] p8 = (((^(5'sd14))?((3'd6)!==(5'd12)):(!(2'd0)))?(&((+(5'sd4))|((5'd23)<<<(4'd11)))):(~|((~(-2'sd1))*(|(4'd6)))));
  localparam signed [3:0] p9 = (~{{((3'd2)<=(3'd4)),(~^(2'd1)),(&(4'd6))},(|(!{{(4'd10),(2'd3),(3'd5)}}))});
  localparam signed [4:0] p10 = (!(3'd4));
  localparam signed [5:0] p11 = (((~^(5'd7))?(+(5'd22)):((2'd0)?(4'd1):(4'd1)))>=(((3'sd2)>>(3'd5))+((4'd13)?(2'd2):(2'd3))));
  localparam [3:0] p12 = (-(4'd2 * (2'd1)));
  localparam [4:0] p13 = ({(2'sd0),(-2'sd0)}?{3{(3'd4)}}:{(4'd7)});
  localparam [5:0] p14 = (({(-4'sd2),(2'sd1)}&{(2'sd0),(2'd2),(5'd19)})|{2{{4{(4'sd1)}}}});
  localparam signed [3:0] p15 = ((((-5'sd1)|(4'd3))>>>((5'sd13)===(5'sd15)))?({4{(2'sd1)}}||((-4'sd0)+(-4'sd2))):(((5'd25)?(3'sd2):(5'd26))=={4{(-5'sd10)}}));
  localparam signed [4:0] p16 = (~({4{((4'sd1)>(3'sd0))}}^~(((4'sd3)>>(-4'sd7))|(4'd2 * (3'd7)))));
  localparam signed [5:0] p17 = (4'd15);

  assign y0 = {4{a0}};
  assign y1 = (~|((+(|(p0^~b1)))<<(~&(-4'sd6))));
  assign y2 = {$unsigned({3{(b1)}}),{(5'd2 * {b2,b2})}};
  assign y3 = ((p6+p6)<(p8?p1:p13));
  assign y4 = ((~^(b0?p15:b1))?(^(~&(b0?a4:b5))):((p5^a2)?(-4'sd6):(a3*b1)));
  assign y5 = (&$signed($signed(((~&a3)+(b4&a0)))));
  assign y6 = {b5,b2};
  assign y7 = (-(3'd1));
  assign y8 = ((~&a4)?(b1<a1):{a1,a1});
  assign y9 = (&p5);
  assign y10 = ((~|(p17+b1))?(p3>a5):({p17,p7}));
  assign y11 = {2{{((b1-b0)!==(~^a5)),{{{b3}}}}}};
  assign y12 = $unsigned((($unsigned(((a1-b3)^~(a3?a1:b2)))===((5'd2 * a0)<<<(a0<=a0)))+($unsigned((p8!=b1))?((p0<=p10)):(p11?p9:p17))));
  assign y13 = {2{(4'd8)}};
  assign y14 = ((((a0?a3:p16)>>>$unsigned(b0))&&(($signed(b0)&&(a1<a2))))>>>(((a2?b4:p11)<(b0?a2:b5))+((a5||b4)!==$signed(b3))));
  assign y15 = (~^(p6?p11:p4));
  assign y16 = (~^(~(~(~|(+(~|(+a3)))))));
  assign y17 = (a1?a2:a5);
endmodule
