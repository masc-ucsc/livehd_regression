module expression_00427(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(&((4'd2)?(+(4'd3)):((2'd0)?(4'sd1):(-2'sd0)))));
  localparam [4:0] p1 = (~^{(!((5'd8)==(5'd26)))});
  localparam [5:0] p2 = (-5'sd3);
  localparam signed [3:0] p3 = ((&(~|(2'sd0)))===(|{4{(4'd0)}}));
  localparam signed [4:0] p4 = {(6'd2 * (3'd4)),(~&(-2'sd0))};
  localparam signed [5:0] p5 = {{(5'sd13),(5'd13)},((5'd10)?(2'd2):(-2'sd0)),(~&(5'd1))};
  localparam [3:0] p6 = ({(-5'sd6)}<((-2'sd1)&(3'd4)));
  localparam [4:0] p7 = ((3'sd2)<<(2'sd1));
  localparam [5:0] p8 = ((((2'sd1)|(2'sd1))||((4'd1)==(4'd9)))===(((5'd31)<=(-4'sd1))>((4'd9)^(-2'sd0))));
  localparam signed [3:0] p9 = ((2'd3)<<<(4'd6));
  localparam signed [4:0] p10 = ((5'd19)==(3'd5));
  localparam signed [5:0] p11 = ((((-3'sd1)<<(5'd30))&(3'd6))===((3'd0)>=((2'd3)<(3'sd2))));
  localparam [3:0] p12 = (-2'sd1);
  localparam [4:0] p13 = {4{({2{(3'd0)}}!=(+(4'sd4)))}};
  localparam [5:0] p14 = (~({(3'd3),(3'sd2),(5'sd1)}>>{(-(2'd2))}));
  localparam signed [3:0] p15 = ((5'd16)*((-3'sd2)?(3'd4):(-5'sd13)));
  localparam signed [4:0] p16 = (~&(((-3'sd1)!==((5'd0)?(3'sd1):(2'd2)))^~((2'sd1)>((3'sd2)?(5'd6):(5'd0)))));
  localparam signed [5:0] p17 = (((-5'sd1)^~(-3'sd3))<<((5'd11)!=(4'sd2)));

  assign y0 = ((~&(((3'd5)|(~&b5))>(-5'sd7)))+(-((b3>b2)?(|(3'd0)):(b0?a3:b5))));
  assign y1 = (-$unsigned((4'd2 * (a2&p2))));
  assign y2 = (~^(~^(+{(a3==a0),{(b0<a4)},(b2|p1)})));
  assign y3 = ((b4?p2:b0)?(p0?a1:p4):{3{p10}});
  assign y4 = (2'd1);
  assign y5 = {1{(((~|{1{a5}})<<<(b0<=b2))+{2{{1{(a5<<p5)}}}})}};
  assign y6 = (+((!(5'd15))+(~(&p10))));
  assign y7 = (5'd2 * (!(b0>>>p8)));
  assign y8 = (~^(~^((-(!(^{4{p4}})))?((p8?a0:a0)>>>(3'd2)):(-4'sd5))));
  assign y9 = (&(~((^(~&(p4>p5)))?((!a4)?{p10,p2,p1}:(!p9)):(&{p6,p10,p8}))));
  assign y10 = (((|(a1^p9))|(p0>>p1))>>(+(2'd2)));
  assign y11 = {1{((~{2{(a0?b2:a0)}})?{4{{b4}}}:(2'd0))}};
  assign y12 = ((p13>p16)?(p6<p15):(a4>=p7));
  assign y13 = (4'd2 * {2{p14}});
  assign y14 = (-4'sd5);
  assign y15 = ((p17?b5:p15)?(3'd0):(3'd1));
  assign y16 = {1{p15}};
  assign y17 = (((~|(2'd0))===(b3>a2))?((a3<=p14)>>>(a2+p5)):((p5<<p6)?(5'sd11):(-p17)));
endmodule
