module expression_00414(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((!((2'sd0)<=(3'd5)))<<<(((-4'sd3)==(5'd8))&&(5'd15)));
  localparam [4:0] p1 = {(~&(-3'sd1))};
  localparam [5:0] p2 = (+(~(|(^((4'sd0)>>>(5'd2))))));
  localparam signed [3:0] p3 = (5'd2 * (&(!(2'd1))));
  localparam signed [4:0] p4 = (~^(^((~&(~(|(4'd15))))!=(+(!(~|(5'sd0)))))));
  localparam signed [5:0] p5 = (-5'sd11);
  localparam [3:0] p6 = (((-2'sd1)/(2'sd1))^(((-5'sd8)^(2'd3))===(!(~&(3'd2)))));
  localparam [4:0] p7 = {4{(-5'sd3)}};
  localparam [5:0] p8 = (~&(4'sd5));
  localparam signed [3:0] p9 = (-((4'd9)?(4'd13):(4'd3)));
  localparam signed [4:0] p10 = ({(3'sd1),(-2'sd0)}?{(4'd14),(2'sd0)}:((5'sd10)>(2'd1)));
  localparam signed [5:0] p11 = {1{{3{((4'd4)||(-4'sd3))}}}};
  localparam [3:0] p12 = {1{(((5'sd12)&&(~((-5'sd13)>(4'd4))))^{3{(&(2'd0))}})}};
  localparam [4:0] p13 = ({((5'd16)==(4'd14))}>=((5'd27)!=(5'd15)));
  localparam [5:0] p14 = ((((4'sd6)|(-3'sd3))>((2'd0)<=(5'sd4)))?({4{(5'd2)}}<{2{(3'sd3)}}):((4'sd7)?(3'd3):(3'd1)));
  localparam signed [3:0] p15 = ({4{(4'd9)}}===(~|{4{(3'sd1)}}));
  localparam signed [4:0] p16 = ((4'd10)!==(((3'd5)===(2'd0))?((-2'sd1)!==(2'd2)):(-4'sd0)));
  localparam signed [5:0] p17 = ((5'd8)?((3'd1)?(-3'sd3):(2'd1)):{(2'd1),(-5'sd15),(5'sd2)});

  assign y0 = ({3{(^(b3<<<p16))}}>=(|{4{$unsigned(p5)}}));
  assign y1 = {{{p2}},{p13,p11,p0}};
  assign y2 = ((-2'sd1)&(~^(4'sd6)));
  assign y3 = {(b3===a2),{a3}};
  assign y4 = (~|{1{{4{{4{p17}}}}}});
  assign y5 = {($unsigned(a0)&$unsigned(b1)),{(a5?b2:b2)},((b0&a0))};
  assign y6 = {4{(~|{p9,p4})}};
  assign y7 = (&{$unsigned((!$unsigned(a5))),((~^{a3})),$unsigned((|(^a5)))});
  assign y8 = {3{{p11,a4}}};
  assign y9 = (-4'sd3);
  assign y10 = ((p12?b2:p17)<<<{1{{1{(-a3)}}}});
  assign y11 = (-((-(~|(+((~&b2)+(+b2)))))===(((!b2)!=(b2-b2))>{(a0+a1)})));
  assign y12 = {($signed({3{p7}})^~(~|(p4?p11:p17))),{4{(p14<<p8)}}};
  assign y13 = {1{(~|{3{$unsigned({b3,a2})}})}};
  assign y14 = (b5+b3);
  assign y15 = (5'd2 * p2);
  assign y16 = ((|(p13&p7))>=(|{b0}));
  assign y17 = (((-4'sd1)===(~^a0))>=((-2'sd0)!==(+b4)));
endmodule
