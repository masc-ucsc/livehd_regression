module expression_00041(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(-5'sd5),(3'sd2),(3'd1)},((5'sd12)||(3'd4)),{2{(3'd4)}}};
  localparam [4:0] p1 = (-(^(!{((-5'sd15)-(-3'sd2))})));
  localparam [5:0] p2 = {4{{2{{1{(4'd5)}}}}}};
  localparam signed [3:0] p3 = ((~|(((-3'sd3)+(2'sd0))>>((5'd13)>>>(4'd3))))==(((4'd1)&(4'sd0))>(^((5'sd5)===(4'd0)))));
  localparam signed [4:0] p4 = {((5'sd6)?(-2'sd0):(3'd5))};
  localparam signed [5:0] p5 = (|(-5'sd6));
  localparam [3:0] p6 = {4{((5'sd13)?(-3'sd3):(3'sd2))}};
  localparam [4:0] p7 = ({2{(4'd14)}}+((4'd1)<<(-3'sd3)));
  localparam [5:0] p8 = ({1{((3'sd3)>=(2'd2))}}>>>((-2'sd0)?(2'd2):(2'd1)));
  localparam signed [3:0] p9 = ((~&{3{(-2'sd1)}})!=(~{2{{3{(-2'sd1)}}}}));
  localparam signed [4:0] p10 = {3{(-3'sd3)}};
  localparam signed [5:0] p11 = {2{{4{(4'sd7)}}}};
  localparam [3:0] p12 = (^({2{{4{(3'd6)}}}}&{4{(5'sd6)}}));
  localparam [4:0] p13 = (~((~(5'sd10))?((-3'sd3)?(2'd2):(3'sd2)):(~|(4'sd1))));
  localparam [5:0] p14 = ({{1{(-4'sd6)}},((4'd13)?(4'sd4):(-4'sd0)),((2'd2)<<(2'd1))}^(((2'd2)-(2'sd0))?((-5'sd7)>>(5'd7)):(-(2'sd0))));
  localparam signed [3:0] p15 = (((2'd2)===(3'd4))^((3'd5)===(4'sd1)));
  localparam signed [4:0] p16 = ({((3'd0)===(2'd1)),{3{(-5'sd4)}}}==(~(((5'd3)||(4'd13))^((2'd1)<(5'd2)))));
  localparam signed [5:0] p17 = (5'sd1);

  assign y0 = (($signed(b0)<(5'sd8))!=$signed((a2?a4:a2)));
  assign y1 = (!(-2'sd1));
  assign y2 = (~^(~((!(a3^~b4))^(^(a5==b1)))));
  assign y3 = ((((p4>>p10)||(p6>p0))^(5'd2 * (b2!==b2)))<({{p5},{p8}}<=({p2}<(p11>b2))));
  assign y4 = {1{(({1{(a3&p0)}}<<(b2^~p13))|{3{(p4^~p17)}})}};
  assign y5 = (~|($unsigned(a3)-(!a2)));
  assign y6 = (((a1?p9:b2)&&(p3?a4:a3))^~((p14<p10)?(p10?b3:p8):{b3,p1}));
  assign y7 = {3{((~&(~^b2))||(~^(^b0)))}};
  assign y8 = {2{{2{{3{p10}}}}}};
  assign y9 = {1{(-{{3{(&{3{b5}})}}})}};
  assign y10 = (-2'sd0);
  assign y11 = (a5?p16:a3);
  assign y12 = (~&(6'd2 * (b2?a2:a1)));
  assign y13 = ((!({$signed(p15)}>>>$unsigned((+a4))))-(((p7-b3))||({p1,p3,p7}==(p16<<b4))));
  assign y14 = ((4'd4)?((p0-p8)&&(p17^~p9)):(p8?p1:p10));
  assign y15 = (2'sd1);
  assign y16 = (-3'sd3);
  assign y17 = ((-(3'd2))-(~((|(b0==a0))-(4'd13))));
endmodule
