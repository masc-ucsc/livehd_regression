module expression_00159(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd0);
  localparam [4:0] p1 = {(-(2'sd0)),(~(2'd3))};
  localparam [5:0] p2 = (|({1{{4{(3'sd2)}}}}<=((3'sd3)?(4'sd5):(-4'sd4))));
  localparam signed [3:0] p3 = (+((!(-(5'd20)))?(-4'sd1):(+((5'd18)>>>(-2'sd1)))));
  localparam signed [4:0] p4 = (-5'sd7);
  localparam signed [5:0] p5 = {3{{4{(4'd11)}}}};
  localparam [3:0] p6 = (!(&((!(&((~(2'd3))&(~^(3'd6)))))>=(~&((~^(5'd26))||((-2'sd0)<=(-4'sd3)))))));
  localparam [4:0] p7 = (&((~&(~|({(-4'sd5),(2'd0),(4'd4)}<(+(-5'sd8)))))+({(-5'sd10),(-5'sd6),(4'd0)}?(-(3'd1)):(+(4'sd3)))));
  localparam [5:0] p8 = {{4{{3{(4'd3)}}}},(3'sd3)};
  localparam signed [3:0] p9 = ((3'sd3)||((5'sd4)&&(-4'sd4)));
  localparam signed [4:0] p10 = {({(5'd31),(3'd4)}-{(2'sd0),(2'd3)}),({(2'd1),(-2'sd1)}||{(-5'sd14),(2'd1),(2'sd1)}),({(-5'sd14)}<{(3'd2),(-4'sd5),(3'sd2)})};
  localparam signed [5:0] p11 = (((3'd3)?(4'd1):(-2'sd0))?((3'd3)&(4'd9)):((-2'sd0)?(3'sd0):(2'd0)));
  localparam [3:0] p12 = (-(((&(5'sd10))&&((-2'sd0)%(3'sd2)))==((-(2'd2))>>>((-3'sd3)!=(3'sd2)))));
  localparam [4:0] p13 = (((-5'sd5)^~(-5'sd15))%(3'd1));
  localparam [5:0] p14 = (5'sd11);
  localparam signed [3:0] p15 = {3{{2{(-4'sd6)}}}};
  localparam signed [4:0] p16 = (~(^(|(~(^(!(^(!(~^(~(-5'sd15)))))))))));
  localparam signed [5:0] p17 = ((5'd25)?(5'd12):(3'd1));

  assign y0 = (((p11>=p16)?(p3?p9:p15):(p15<<b5))>>$unsigned(($signed($signed((a2!==a2)))|($unsigned($signed(a0))))));
  assign y1 = (-b1);
  assign y2 = (((2'd0)?(a4+a1):(~^p9))^~((p3==p14)?{p2,a3}:(~p6)));
  assign y3 = (((-{3{a5}})?{1{(a4||p8)}}:(&{4{p14}}))-{1{(~{4{(b3?a3:a1)}})}});
  assign y4 = {2{({a0,p1}>={4{p13}})}};
  assign y5 = ((^p17)?(p9^p0):(!p11));
  assign y6 = ((p6?a1:p9)?((b2!==b1)&(b0?p7:p6)):(a1?p15:p0));
  assign y7 = {(p2|p7),{2{p8}}};
  assign y8 = ($unsigned((((3'sd3)===(!a3))||$signed((^(b2<a1)))))&&{3{(a1==p12)}});
  assign y9 = (-((~|b5)&&(&b3)));
  assign y10 = (3'sd1);
  assign y11 = (4'd6);
  assign y12 = ({4{{4{a0}}}}?((p15>p2)^~(p3||b0)):(~&((b2!=a5)>=(b1>>a0))));
  assign y13 = ({1{((b4?b4:a5)?(b1===a1):{1{{4{b2}}}})}}>{1{((b4?b1:b0)+({2{a0}}>>>(b0>>b1)))}});
  assign y14 = {(^(!{{{{b0,p9},{a0}},{p16,p14,p2}},(~^{{p14,p13,b0},(&a2),{b4,p2}})}))};
  assign y15 = (~&(+$unsigned((-5'sd15))));
  assign y16 = (6'd2 * b0);
  assign y17 = $unsigned((^((p11==p14)^(^(4'd4)))));
endmodule
