module expression_00753(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~^(^((-5'sd13)?(4'd3):(-2'sd0))))?(-(&((3'sd0)>>(4'd13)))):((3'd0)?(5'd21):(2'd2)));
  localparam [4:0] p1 = (|(((-4'sd1)?(5'd24):(3'd2))/(5'd4)));
  localparam [5:0] p2 = (!(^((4'sd4)&&(-2'sd0))));
  localparam signed [3:0] p3 = (((3'd2)?(3'd7):(4'sd2))!=(~((4'd12)<<(3'd0))));
  localparam signed [4:0] p4 = {3{((3'd1)<=(4'd11))}};
  localparam signed [5:0] p5 = {{{4{((-5'sd4)?(3'd5):(-3'sd1))}}},(2'd3)};
  localparam [3:0] p6 = {3{(|(~{4{(5'sd6)}}))}};
  localparam [4:0] p7 = (~|(^((^{((3'd1)!==(3'd3))})>(!{{3{(-2'sd1)}}}))));
  localparam [5:0] p8 = (|(((+((3'd5)!=(2'sd0)))!=((4'd9)?(4'd0):(-3'sd1)))|(((5'sd8)-(4'sd0))<<(~(~|(2'd2))))));
  localparam signed [3:0] p9 = (5'd2 * ((2'd2)?(2'd3):(3'd1)));
  localparam signed [4:0] p10 = ((^(-{({(5'sd12),(3'sd0),(2'd3)}==={(-4'sd7),(-3'sd0),(4'd4)})}))<<<(~{((5'd2)-(-2'sd0)),(&(3'sd0)),{(4'sd5),(2'd1),(-3'sd2)}}));
  localparam signed [5:0] p11 = (5'sd5);
  localparam [3:0] p12 = ((+(3'd7))!=={2{((-3'sd3)<<<(-3'sd0))}});
  localparam [4:0] p13 = {4{(5'sd12)}};
  localparam [5:0] p14 = {2{{{4{(-2'sd0)}},{(2'd3),(4'sd0)},((-5'sd10)>>(5'd19))}}};
  localparam signed [3:0] p15 = ((((2'd0)||(5'sd3))==((3'd4)&(-2'sd0)))-(((5'd9)<<<(5'd20))<<<((4'd1)%(3'd4))));
  localparam signed [4:0] p16 = ({(5'd18),(5'sd11),(-5'sd1)}?{(2'd1),(5'd14),(5'sd14)}:(((5'sd15)?(3'd6):(-2'sd1))!==((4'sd2)>=(2'd0))));
  localparam signed [5:0] p17 = (&(-(~&(((&(2'sd0))<((-4'sd3)^(-4'sd5)))<<(~|((3'd6)*(4'd6)))))));

  assign y0 = (((b0^~b2)&(a1>=a2))<<{((b3?b0:a3)>>{b4,b5})});
  assign y1 = (+((a0^p16)==(~p9)));
  assign y2 = (6'd2 * (a0+p1));
  assign y3 = (-(-5'sd10));
  assign y4 = {3{{3{p7}}}};
  assign y5 = (&((4'sd6)^~(p8&p6)));
  assign y6 = {2{(+(6'd2 * p6))}};
  assign y7 = (&(a0?a2:b2));
  assign y8 = (5'sd7);
  assign y9 = (((p1&p5)<=(&p10))?((a0||p1)>{4{p4}}):(^(-(a2===a5))));
  assign y10 = (~^(~&{a0,b3,p14}));
  assign y11 = $unsigned(({2{(&{3{p10}})}}?((~(-2'sd0))):({1{p1}}?(p3?p6:p16):(p10))));
  assign y12 = ((~&b5)&&(~^p12));
  assign y13 = {3{b4}};
  assign y14 = {{{(a1>b2),(!p4),(~p5)},((^(!a3))===({a5})),((-(|$signed((|(-p13))))))}};
  assign y15 = (5'd21);
  assign y16 = {b3,b4};
  assign y17 = ({1{a4}}!==(5'd2 * b0));
endmodule
