module expression_00796(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((((2'd0)!==(-4'sd3))^((3'sd1)==(3'd4)))?(((4'sd2)?(2'd0):(3'd0))?{3{(3'd1)}}:((-2'sd0)>>(4'd5))):(((2'd1)>>>(2'sd0))=={(5'sd9),(4'd11)}))};
  localparam [4:0] p1 = (((2'sd1)!=(2'd2))==((3'sd3)!=(3'd4)));
  localparam [5:0] p2 = (!(2'd2));
  localparam signed [3:0] p3 = ((((5'd31)===(-4'sd2))>>>((3'sd1)?(3'sd3):(5'sd3)))>>(~|((5'd11)<=(4'd5))));
  localparam signed [4:0] p4 = (~(5'sd15));
  localparam signed [5:0] p5 = {1{{4{(2'd0)}}}};
  localparam [3:0] p6 = (~|(2'sd1));
  localparam [4:0] p7 = (~&(5'd3));
  localparam [5:0] p8 = (~(~|(2'd3)));
  localparam signed [3:0] p9 = {(-4'sd7),(5'd30)};
  localparam signed [4:0] p10 = ((+(((3'sd1)<(4'sd5))?((4'd9)||(-2'sd0)):(^(4'sd4))))===(((5'd30)?(2'd1):(5'd28))&&(((2'd2)<<<(4'd4))&&((2'sd0)<<(5'd29)))));
  localparam signed [5:0] p11 = (-(~(3'd5)));
  localparam [3:0] p12 = (+(((+(^(3'd1)))/(4'sd5))&(((-5'sd14)<<(-5'sd7))!==(!((-3'sd2)>>(3'd0))))));
  localparam [4:0] p13 = (~&(^((((3'd3)<<(3'd4))>(+(~(3'd0))))<=(((-2'sd0)&(2'd1))-(!(~(3'sd1)))))));
  localparam [5:0] p14 = {4{(~&(3'd3))}};
  localparam signed [3:0] p15 = {1{(({3{(4'd1)}}<<<((-3'sd1)!=(3'd2)))&&(4'd2 * ((2'd3)+(5'd25))))}};
  localparam signed [4:0] p16 = (6'd2 * ((3'd1)?(4'd4):(2'd3)));
  localparam signed [5:0] p17 = {4{(5'd7)}};

  assign y0 = ((~&(a2>>b0))===(a4-b3));
  assign y1 = (~^((a1&p10)/a0));
  assign y2 = (|{4{(!($signed(p12)))}});
  assign y3 = $unsigned(({{p4,p14,a4},(a5!==a3),$unsigned((p7))}|($unsigned((p9|p4))&((a3|p0)))));
  assign y4 = (((~&a1)?(^p5):{1{a1}})?(~^(~{2{(~^b3)}})):({2{a3}}?(|a2):(p1?b0:b0)));
  assign y5 = ((-(~(2'd1)))<(-(~(a0!==a0))));
  assign y6 = (~^(+(~(~(&(|(~(|(~^(3'sd1))))))))));
  assign y7 = ((+((p0<<<p8)||(p10?b0:a4)))?((b5/b4)/p13):($signed(b5)&&(~p11)));
  assign y8 = (6'd2 * (p2?b1:b2));
  assign y9 = {4{(~|$unsigned((!b4)))}};
  assign y10 = {4{(-3'sd1)}};
  assign y11 = (({2{b0}}?(b1>>p17):(4'sd6))>((a4?b3:a2)?{2{b0}}:(b3>b0)));
  assign y12 = {{4{p16}},((~a4)<<<{2{p7}})};
  assign y13 = (2'd1);
  assign y14 = ((p4%p9)-$unsigned((p13)));
  assign y15 = ((p4?b5:b2)?(~^b0):{2{p17}});
  assign y16 = ((a0>>a2)!==(a5&&a3));
  assign y17 = ((4'd2 * (a1?p8:p13))?{b2,a4,a3}:(+(~&{p2})));
endmodule
