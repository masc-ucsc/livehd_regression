module expression_00533(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd1);
  localparam [4:0] p1 = {4{{2{(4'sd2)}}}};
  localparam [5:0] p2 = ((5'd10)>=(-5'sd3));
  localparam signed [3:0] p3 = (~&((6'd2 * (4'd9))<<(-((2'd3)?(3'd6):(3'd3)))));
  localparam signed [4:0] p4 = {1{(((2'd2)?(-5'sd11):(4'd9))?{4{(5'sd4)}}:{4{(5'd16)}})}};
  localparam signed [5:0] p5 = ((+(5'd8))^(~|(-3'sd0)));
  localparam [3:0] p6 = ({((&{(4'd4),(5'd1)})===(&((-5'sd0)^(3'd1))))}<={(3'd5),((2'sd0)<=(4'sd2))});
  localparam [4:0] p7 = (-(~&(((~&(4'd3))!=((-2'sd0)||(3'd4)))<((~&(3'd4))===(|(3'd4))))));
  localparam [5:0] p8 = (3'd2);
  localparam signed [3:0] p9 = {4{(-4'sd4)}};
  localparam signed [4:0] p10 = {{(!{(3'd5)}),(&(&{{(2'sd0),(5'd11),(4'd1)}})),(~(+{(-3'sd0),(4'sd4),(5'd27)}))}};
  localparam signed [5:0] p11 = (((5'd5)-(|(5'd6)))^~((+(5'd0))!==((3'd2)&(2'd0))));
  localparam [3:0] p12 = (|(3'd6));
  localparam [4:0] p13 = {4{(4'sd7)}};
  localparam [5:0] p14 = {(-5'sd2),(-3'sd3),(2'd0)};
  localparam signed [3:0] p15 = (~&{1{{4{(5'd18)}}}});
  localparam signed [4:0] p16 = ({(6'd2 * (5'd6)),{4{(4'd6)}}}===(((2'sd1)==(4'd1))=={4{(2'd0)}}));
  localparam signed [5:0] p17 = (!(3'd6));

  assign y0 = (!{3{(2'sd0)}});
  assign y1 = (((b5>>a1)?(b1<<b5):(a5?p0:a0))>>>((5'sd15)<=(-5'sd12)));
  assign y2 = ($signed(($unsigned((|{(p4==p1),(~|{p13,a5,p12})}))^~($unsigned({p10,b3,b5})>>>{{p14},{p9,p5,p4}}))));
  assign y3 = ((5'd2 * (b2!==b2))<(((b2&a5)^(a1?p4:b5))|((b2<<b3)^~(b5%a0))));
  assign y4 = (~&{(+p12),(!p2)});
  assign y5 = (((p3?p15:p17)?{p6,p12}:(p12?p4:p4))?({4{p10}}?{4{p10}}:{p5}):{4{p16}});
  assign y6 = {4{($signed(p8)>>>(^b4))}};
  assign y7 = {4{(a4?a0:a0)}};
  assign y8 = (~(((^{1{(|(p16^p3))}})>=((2'd2)!==(b2>>>a2)))!=(((2'd2)<{p16,p5})^~(5'd22))));
  assign y9 = {1{((2'd3)&&(-3'sd2))}};
  assign y10 = ({{b5,b1},(!{b5,p0,b0})}?{$unsigned((^(a2?a1:b1)))}:$signed((~^(~$unsigned((-(&a3)))))));
  assign y11 = {{3{(a1>>>a2)}}};
  assign y12 = (!$unsigned((&$signed((-4'sd0)))));
  assign y13 = (~^(~(~&(b2^~b5))));
  assign y14 = (({3{b3}}^~((a4&&a1)==={a4,a0,b5}))<<<(({p3,a5}||{p13,p1,a0})||{4{p10}}));
  assign y15 = ((b3>p11)||(b1>=a1));
  assign y16 = (~&(p11>>>p1));
  assign y17 = {b5,a5};
endmodule
