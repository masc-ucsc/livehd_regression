module expression_00968(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((2'd2)+(-2'sd1))||((5'd2)===(3'd1))),{(^((3'sd1)-(-2'sd0)))},(~^((~(4'sd0))>=((2'd0)>>(3'sd2))))};
  localparam [4:0] p1 = ((2'd0)>=(3'd1));
  localparam [5:0] p2 = (~^(({(5'sd3),(-3'sd0)}&&{(4'sd5)})==((&(-3'sd0))>>>(4'd15))));
  localparam signed [3:0] p3 = {4{(-2'sd0)}};
  localparam signed [4:0] p4 = (2'd3);
  localparam signed [5:0] p5 = (^((5'd2 * (3'd7))>>((-4'sd6)==(-5'sd12))));
  localparam [3:0] p6 = ((-4'sd0)?(2'd0):(4'd5));
  localparam [4:0] p7 = {(2'd2)};
  localparam [5:0] p8 = {((~&(2'd3))?(~^(5'd8)):{(4'sd6)}),((-(2'sd1))?(^(2'd1)):{(2'd3)}),({(-3'sd2)}?{(2'sd1),(3'd6),(2'sd1)}:((5'd18)?(5'sd15):(3'd1)))};
  localparam signed [3:0] p9 = (((4'd9)>(3'd6))?((5'sd4)?(5'sd8):(5'd29)):(|((-4'sd3)&(3'sd2))));
  localparam signed [4:0] p10 = (((3'd1)===(2'd0))<=((5'sd3)<(-3'sd1)));
  localparam signed [5:0] p11 = {3{(-(5'd3))}};
  localparam [3:0] p12 = {{(2'sd0),(3'sd2),(2'sd1)}};
  localparam [4:0] p13 = (-{(&(3'sd3))});
  localparam [5:0] p14 = {({3{(2'd2)}}!=={(5'sd2),(3'd7),(4'd15)}),{2{(-5'sd3)}},(3'sd2)};
  localparam signed [3:0] p15 = (((4'd8)?(-3'sd2):(-2'sd0))+{4{(4'd1)}});
  localparam signed [4:0] p16 = {({((5'd30)&(-3'sd3)),((2'd1)?(-4'sd6):(5'd6))}<<<({(5'd24),(3'd4),(4'sd7)}?((-3'sd1)?(2'sd1):(2'd3)):((2'sd0)===(3'd7))))};
  localparam signed [5:0] p17 = {(4'sd5),(4'd2),(-5'sd5)};

  assign y0 = {2{{(-3'sd1),(a4^p9),(3'd0)}}};
  assign y1 = (5'd19);
  assign y2 = $signed((~|(p11^p17)));
  assign y3 = (b4|a3);
  assign y4 = ((-p13)?(b1?a4:b3):(-a3));
  assign y5 = ((3'd1)?(~^(a3?p13:a5)):(~&(p3?a0:a0)));
  assign y6 = ({2{{4{p16}}}}-({2{p11}}>>>{p5}));
  assign y7 = {{1{{1{{(|{1{(!(~&{p11,a2,b3}))}}),(!(^{(~b2),{a3,p1,a5}}))}}}}}};
  assign y8 = ({4{p17}}<(p5>p8));
  assign y9 = (((~&(p0&p2))==($unsigned(p11)<<<{4{p10}}))&&((^(~|{1{p15}}))+($signed(p1)=={1{p16}})));
  assign y10 = {1{(p1||a4)}};
  assign y11 = (((|b2)<<(|p3))^(!{2{(|p15)}}));
  assign y12 = (~&{((-(~p2))>>(+(a0<<<p3))),(~&(((+b2))!=={b0,b1}))});
  assign y13 = $unsigned((2'd0));
  assign y14 = (((b4?b3:a3)?(a4?a2:p5):(p5?b5:b2))==((p12>>>p6)?(b5?a0:b0):(a4?p1:a3)));
  assign y15 = (((-a2)));
  assign y16 = (-3'sd0);
  assign y17 = {2{{3{(~^(~&p11))}}}};
endmodule
