module expression_00823(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(~|(|(^(+(2'sd1))))));
  localparam [4:0] p1 = ({{(4'd10),(3'd1)},((3'sd3)<(5'd25)),((5'sd6)<=(2'sd1))}<=({(2'd1),(-3'sd3),(3'd4)}>>((5'd24)<(-2'sd1))));
  localparam [5:0] p2 = (({4{(4'd8)}}^((5'd22)?(-2'sd0):(-5'sd3)))?{2{(~^(5'd13))}}:(|((4'd9)?(-4'sd5):(4'd9))));
  localparam signed [3:0] p3 = {4{((2'sd1)?(4'd8):(4'sd1))}};
  localparam signed [4:0] p4 = ((2'd0)!=={4{(-3'sd0)}});
  localparam signed [5:0] p5 = (+(!(~|(4'sd3))));
  localparam [3:0] p6 = ((((4'd6)!=(-4'sd3))>>((4'd2)?(4'd5):(-5'sd3)))?{4{(5'd24)}}:{{2{{3{(3'd4)}}}}});
  localparam [4:0] p7 = (~&{{3{{4{(2'd3)}}}},(~&{2{((4'd0)?(4'd4):(-3'sd2))}})});
  localparam [5:0] p8 = {3{(4'd15)}};
  localparam signed [3:0] p9 = (5'd2 * ((3'd1)<(3'd1)));
  localparam signed [4:0] p10 = (((~&(2'd3))<=((-3'sd3)?(4'd0):(-5'sd15)))?(+{(2'd0),(-4'sd2)}):{1{((-3'sd0)<=(-4'sd0))}});
  localparam signed [5:0] p11 = ((((5'd13)?(3'd6):(-4'sd1))===((-3'sd1)!==(2'sd0)))<<<(~|(-(4'd2 * ((2'd1)<<(2'd3))))));
  localparam [3:0] p12 = (4'd7);
  localparam [4:0] p13 = (^(5'd25));
  localparam [5:0] p14 = {((-5'sd8)>>(5'd7))};
  localparam signed [3:0] p15 = ({1{((4'd2 * (3'd0))&&((5'sd0)<<(5'sd9)))}}>{3{((-3'sd2)!==(-2'sd0))}});
  localparam signed [4:0] p16 = {3{(2'd3)}};
  localparam signed [5:0] p17 = {2{{2{(~&((-5'sd10)<=(-5'sd14)))}}}};

  assign y0 = (p6?p2:p9);
  assign y1 = (!{a4,a4});
  assign y2 = {$signed((5'sd12)),(^(~|(~{(+p6),(~|a3)}))),$signed({(+b2),(3'sd0),(3'd7)})};
  assign y3 = {4{{1{((p11>>p5)+(p4>>>p8))}}}};
  assign y4 = (-((~&((a4>a3)))|({4{a4}}<(|b2))));
  assign y5 = (~&(((~&p14)||(5'd2 * p12))?(~|(^(~|p14))):(~^(+(~^p6)))));
  assign y6 = (b1<p3);
  assign y7 = $unsigned((|({4{p0}}>>>{3{a5}})));
  assign y8 = {{(p4>p8),(a1<p1)},({p2,p17,a3}==(p5>=a1))};
  assign y9 = {3{(3'd6)}};
  assign y10 = ((-{(^a1),(2'sd0),(!p8)})+(~^(!{a4,b3,a4})));
  assign y11 = (5'd2 * $unsigned((a1<<p5)));
  assign y12 = ({((({p14,p1,p3}>=(p16>>p16))))}&&({a4,b5,a5}===($signed(b4)=={a1,b2,b4})));
  assign y13 = (b3>>>p6);
  assign y14 = (|(~{2{(b5!==b3)}}));
  assign y15 = ({2{p1}}-{4{p9}});
  assign y16 = (~^$unsigned($unsigned(p11)));
  assign y17 = (-4'sd5);
endmodule
