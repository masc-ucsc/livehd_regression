module expression_00301(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{2{(2'd0)}});
  localparam [4:0] p1 = {4{(&((3'd2)<<(3'sd1)))}};
  localparam [5:0] p2 = (((3'd4)?(2'd3):(-2'sd0))>=(~&{3{(3'd5)}}));
  localparam signed [3:0] p3 = ((2'sd1)-(-4'sd1));
  localparam signed [4:0] p4 = (+(^({3{(4'd15)}}===(((2'sd0)<=(4'd0))+{1{(5'sd11)}}))));
  localparam signed [5:0] p5 = (~^((-3'sd3)?(2'd0):(4'sd0)));
  localparam [3:0] p6 = ((4'd4)^(3'sd0));
  localparam [4:0] p7 = {(+{(|(~&(-5'sd3))),(^((-5'sd5)!==(5'd16)))}),((-4'sd7)<(~|(~(&(2'd0)))))};
  localparam [5:0] p8 = (2'sd1);
  localparam signed [3:0] p9 = (-4'sd1);
  localparam signed [4:0] p10 = (5'sd13);
  localparam signed [5:0] p11 = {{1{{3{(5'd13)}}}},{1{(~^(|(2'sd0)))}}};
  localparam [3:0] p12 = ({4{{4{(4'd11)}}}}>>>{4{(^(2'd3))}});
  localparam [4:0] p13 = {{(-4'sd7),(5'sd4)},(~|(-3'sd2))};
  localparam [5:0] p14 = (5'sd8);
  localparam signed [3:0] p15 = ({{(2'd1),(3'd5)},(|{4{(2'd0)}}),{(3'sd3),(5'sd10),(-3'sd2)}}>>(|{1{{4{{3{(4'd9)}}}}}}));
  localparam signed [4:0] p16 = (-4'sd3);
  localparam signed [5:0] p17 = (2'sd1);

  assign y0 = (p6&p8);
  assign y1 = {{$unsigned({p8}),(p3?p1:p13),(p14+p8)},{({p8}<<<(4'd2 * p7)),((p5-p12)&&(p6>>p1))}};
  assign y2 = (~^b5);
  assign y3 = ((-5'sd15)>>(5'd2 * p1));
  assign y4 = $unsigned(((3'sd3)<(((~&(4'd2 * a0)))!==((2'sd0)==(a5!=b3)))));
  assign y5 = (-b0);
  assign y6 = {1{{2{{2{(&(3'sd3))}}}}}};
  assign y7 = (~&(-(~|p7)));
  assign y8 = (~^(~(~(~|(^a5)))));
  assign y9 = ((-3'sd3)-((~&(&{a1}))^~((~|p16)>>>{p7,p12})));
  assign y10 = $unsigned($unsigned($signed((($signed(a2)&&(a4<a4))>>{4{a1}}))));
  assign y11 = (a0?b3:a2);
  assign y12 = (((6'd2 * (p2?p13:p13))&&((p1?p1:a4)>(p9-p7)))^(+((p5&&p5)?(!b2):(p2?p10:a4))));
  assign y13 = (&(((b5>>>p3)/a2)-(^((^b0)||(p2>>>p10)))));
  assign y14 = $unsigned({1{((((~^{4{b2}})>={3{a2}})||($signed((-(b3>>b4)))>>({3{b2}}&(p5<a2)))))}});
  assign y15 = {$signed((5'd30))};
  assign y16 = ((~|(-((a4<p7)>>>(5'sd11))))<<<(&{2{{2{p1}}}}));
  assign y17 = (-3'sd3);
endmodule
