module expression_00425(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd2 * ((4'd8)!=(4'd1)))?(((3'd3)&&(-5'sd12))*((3'd6)+(5'd0))):(((5'd10)/(3'sd0))==((3'sd1)/(2'd2))));
  localparam [4:0] p1 = (((2'd3)?((5'sd11)?(4'sd6):(2'd2)):(&(2'd2)))<<<(((4'd7)?(5'd11):(3'd4))===((4'sd4)===(-5'sd1))));
  localparam [5:0] p2 = ((|(+{{(4'd11),(4'sd7)},(~^(4'd4))}))>=((^{(3'd1),(5'd1)})&{(2'd1),(5'sd14)}));
  localparam signed [3:0] p3 = (4'd0);
  localparam signed [4:0] p4 = (^(5'd5));
  localparam signed [5:0] p5 = ((&(2'd0))^~(-(5'd18)));
  localparam [3:0] p6 = ((-3'sd1)!=(3'sd2));
  localparam [4:0] p7 = {((5'd7)+(5'sd12)),((4'sd2)+(-3'sd3))};
  localparam [5:0] p8 = (6'd2 * ((2'd2)===(2'd1)));
  localparam signed [3:0] p9 = {({(3'd2),(2'sd1),(2'd3)}>>{(5'sd5),(3'd2)})};
  localparam signed [4:0] p10 = {2{((2'd2)<<<(5'd27))}};
  localparam signed [5:0] p11 = (!(~({((4'd14)<<(2'd3))}&{(2'd0),(-3'sd0),(3'd6)})));
  localparam [3:0] p12 = (~^((~^(4'd9))==(3'd7)));
  localparam [4:0] p13 = ((3'd6)<=(-3'sd1));
  localparam [5:0] p14 = ({4{(5'd25)}}?(~(((5'd3)>(4'd9))===((4'd3)?(2'd0):(4'd7)))):{2{((5'd26)?(4'd4):(2'd3))}});
  localparam signed [3:0] p15 = (~^(~^(3'd7)));
  localparam signed [4:0] p16 = (~&{3{(2'd3)}});
  localparam signed [5:0] p17 = ((((5'sd13)||(5'd7))!=(2'sd1))-(((5'd14)===(4'sd0))>>((2'd1)^(5'd13))));

  assign y0 = ((b1?a1:a4)>>>(a3>=b3));
  assign y1 = (|({(b3<<a4),(4'sd6)}-(5'd17)));
  assign y2 = (6'd2 * (p12-p8));
  assign y3 = ((a1?p15:b2)?({2{b2}}):(a1==p7));
  assign y4 = $unsigned((((p17?b2:p10)?$unsigned({p4}):{1{(p0<<p1)}})=={1{({3{$unsigned($unsigned(p11))}})}}));
  assign y5 = (({3{b0}}>>>(~&(b1>b4))));
  assign y6 = (^{(~|(p12?p7:p17)),(~|{p11,p2}),(-(a4?p7:p15))});
  assign y7 = ((b0!==a3)<=(-(~|b1)));
  assign y8 = {{b5,p14},{2{a1}},{1{(p10>p17)}}};
  assign y9 = {3{{a3,a0,a0}}};
  assign y10 = {1{({3{{3{b3}}}}==(((-2'sd1)>>{a4})!={(4'd9)}))}};
  assign y11 = ((!((|b5)&&{p0}))?(~|(|(a2?p9:p12))):{(p14>p14),(^p14)});
  assign y12 = (+(^(2'sd0)));
  assign y13 = (~|((b3<<p16)/p4));
  assign y14 = (((!b5)^(a4<=p14))>(&((p4<<p17)<(p13|a4))));
  assign y15 = {3{{p5,p7,p12}}};
  assign y16 = ((~&((b1?b4:p11)?(b3?a0:a3):(b3<=a2)))?((a0||b0)?(|p6):(a1<<<b0)):(~^((a0/a0)?(a5?p4:p14):(~|a5))));
  assign y17 = ((6'd2 * (3'd3)));
endmodule
