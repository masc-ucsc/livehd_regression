module expression_00641(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(4'sd3),(-5'sd1)}>=(~|{(5'd17)}));
  localparam [4:0] p1 = (-((-(((5'sd10)!=(4'd9))-((4'd11)<<(4'd7))))==(3'd1)));
  localparam [5:0] p2 = (((&(3'sd1))>(4'd15))||(~&(^((-4'sd0)!=(3'sd3)))));
  localparam signed [3:0] p3 = (+((&{(-4'sd1),(3'sd2),(3'd6)})>>>(3'd3)));
  localparam signed [4:0] p4 = {(({(-3'sd0),(4'd2),(3'd0)}?((-5'sd8)<<<(2'sd0)):(5'd2 * (2'd1)))?({(3'd0)}<((3'd1)<<<(2'd0))):{{(5'd24),(5'd25)},((2'd1)?(5'd8):(-2'sd0)),(+(5'd3))})};
  localparam signed [5:0] p5 = (~(-3'sd2));
  localparam [3:0] p6 = (~|(((4'sd1)?(5'd25):(-5'sd11))?(~&{3{(4'd13)}}):(^((-4'sd5)-(2'd1)))));
  localparam [4:0] p7 = (3'd2);
  localparam [5:0] p8 = ((6'd2 * ((5'd31)>=(3'd4)))=={1{(((2'sd1)<(3'd5))!=((5'sd1)^(-5'sd2)))}});
  localparam signed [3:0] p9 = (~{2{{4{(~^(2'sd1))}}}});
  localparam signed [4:0] p10 = ((4'sd0)?(3'd3):(5'd13));
  localparam signed [5:0] p11 = (((3'd1)===(2'd1))|(&((5'd21)>>(2'd2))));
  localparam [3:0] p12 = {3{{3{(3'd0)}}}};
  localparam [4:0] p13 = (2'd1);
  localparam [5:0] p14 = (((5'd28)&((5'd10)&(-2'sd1)))<=(~|{((3'd3)+(-4'sd3)),(-4'sd7),((-4'sd4)>>(-2'sd1))}));
  localparam signed [3:0] p15 = (+({3{(~(3'd6))}}?(~^(~&{1{(4'd2 * (2'd0))}})):(((4'd11)<<<(4'd10))<(5'd2 * (5'd9)))));
  localparam signed [4:0] p16 = ((~&(|((3'd3)&(5'd28))))^(((-4'sd0)%(-5'sd7))<=((5'd14)-(2'd2))));
  localparam signed [5:0] p17 = (-4'sd0);

  assign y0 = ((((a4!=b1)===(b2>>b4))!==((a0==a2)>>(a2>>>b0)))^~(((p2<<b0)+(b1===b4))&&((a2||b2)!==(b4||b0))));
  assign y1 = (|(5'd5));
  assign y2 = (((a1&&a0)||(b4||b3))!==$unsigned((-2'sd0)));
  assign y3 = (((~(^b2))&&(~^(b1>>>b1)))===((a3>>>a3)!==(a3&b0)));
  assign y4 = {(5'd27)};
  assign y5 = ((&$unsigned((!(p16&&b4))))?(4'd6):$unsigned((2'sd1)));
  assign y6 = ((a1<<<b2)?(p16?a3:p8):{(a3?p6:a0)});
  assign y7 = (-4'sd4);
  assign y8 = (3'd0);
  assign y9 = (p8?p11:b1);
  assign y10 = (p9&p12);
  assign y11 = ((~|a4)>>{3{b5}});
  assign y12 = (~&(!(~{2{(~(&p10))}})));
  assign y13 = {1{(({4{p16}}<={3{p13}})?({b0}?(p0>>b0):(p6)):((p15?p8:b1)?(b5!==b2):(p17?p2:a0)))}};
  assign y14 = ({a4,p3,b0}&(b4>=p17));
  assign y15 = (((p12?p3:a4)|(-p17))<=((p7^b4)!=(p1>p10)));
  assign y16 = $unsigned({$signed((a1)),$unsigned((p0)),{3{b2}}});
  assign y17 = (!(((~^($unsigned((b1<=p17))+(!(+a0)))))&(&(~|$unsigned((&(~^(!(5'd2 * p8)))))))));
endmodule
