module expression_00711(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{({2{(3'sd2)}}<<((-3'sd1)?(-3'sd3):(3'd2)))}}?(((-4'sd5)>>(3'd3))<{4{(5'd0)}}):(((4'd4)^(-4'sd0))?((-2'sd1)>>(3'd5)):((-3'sd1)?(-2'sd1):(2'sd0))));
  localparam [4:0] p1 = (((+(2'd0))|((2'd0)?(4'sd2):(4'd6)))?({3{(-5'sd8)}}-((3'sd1)>=(3'd0))):({2{(5'sd10)}}>(|(5'd16))));
  localparam [5:0] p2 = ({(4'd7),(4'sd2)}?{((-2'sd1)&(3'd5))}:{4{(3'sd3)}});
  localparam signed [3:0] p3 = {3{({(-5'sd7),(3'd0),(2'd3)}>(4'd2 * (4'd10)))}};
  localparam signed [4:0] p4 = ((5'd1)===(-4'sd6));
  localparam signed [5:0] p5 = (4'd10);
  localparam [3:0] p6 = (5'sd3);
  localparam [4:0] p7 = ({(2'd1),(4'sd7)}<(!((2'd2)?(-4'sd6):(5'sd2))));
  localparam [5:0] p8 = (3'd2);
  localparam signed [3:0] p9 = (5'd13);
  localparam signed [4:0] p10 = {3{((-3'sd1)<=(-2'sd1))}};
  localparam signed [5:0] p11 = ({3{(-5'sd6)}}!==((-2'sd1)&&(-3'sd1)));
  localparam [3:0] p12 = {3{((2'd1)>(4'd12))}};
  localparam [4:0] p13 = {1{({3{{2{(-4'sd1)}}}}&((+{4{(3'd6)}})-{1{((-3'sd1)&(2'd3))}}))}};
  localparam [5:0] p14 = {1{{3{((3'sd0)<<(3'sd3))}}}};
  localparam signed [3:0] p15 = (^({1{((4'sd4)-(3'sd0))}}<<<(-(^((-2'sd1)<<<(5'sd9))))));
  localparam signed [4:0] p16 = ({{3{((3'd6)<=(-2'sd0))}}}&((!(-3'sd2))?((5'd25)<<(3'd6)):(2'd0)));
  localparam signed [5:0] p17 = (^((5'sd14)?(-2'sd0):(3'd5)));

  assign y0 = (~^(3'sd1));
  assign y1 = (((3'sd0)&&(p14<=p0))?((3'sd1)!=(2'sd0)):(-5'sd10));
  assign y2 = ((~&(((~|p15)-(!p15))==(+(p3+p16))))==(!(|($signed((p12|p3))>=(~(p14^p11))))));
  assign y3 = ((((|b5)<={4{a3}})>>((+p11)||$unsigned(p12)))>>(&(!(-($unsigned({2{b3}}))))));
  assign y4 = (~&(-$unsigned(((~&$unsigned((~(|p16))))))));
  assign y5 = (-(+{4{{4{a5}}}}));
  assign y6 = (2'sd0);
  assign y7 = (4'd1);
  assign y8 = (5'd15);
  assign y9 = (((|{2{b4}})&&((!a3)))?({1{{b2,p4}}}&(b4?a2:a0)):(({b4,p14,b0}<={4{p15}})));
  assign y10 = ({3{(3'd2)}}?$unsigned($unsigned({3{p0}})):{4{p0}});
  assign y11 = $signed($signed(($unsigned((~((a4|b3)!==(3'd2))))>(3'sd1))));
  assign y12 = (p1?p12:p0);
  assign y13 = (~^b1);
  assign y14 = (((p8>b0)<(p16|b5))>>($signed((b3&a3))===(~^(~b3))));
  assign y15 = (($unsigned((4'd6))?(a4?p11:b4):(5'sd1))||(3'd7));
  assign y16 = $unsigned((5'd2 * (b0&&p6)));
  assign y17 = ((3'sd3)===(a4+b3));
endmodule
