module expression_00629(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(|{3{{3{(-3'sd1)}}}}));
  localparam [4:0] p1 = (((3'd1)?(5'sd2):(-2'sd1))?((-2'sd1)>=(4'd0)):((2'd3)?(-5'sd9):(4'd3)));
  localparam [5:0] p2 = ((-4'sd2)-(3'sd0));
  localparam signed [3:0] p3 = (-((|(5'sd8))==(!(!((~&(5'd2))|(5'd30))))));
  localparam signed [4:0] p4 = (((-2'sd1)<=(4'd12))*((4'd12)-(-2'sd1)));
  localparam signed [5:0] p5 = (-({2{((-4'sd6)>>(4'd5))}}>>>(|((~&(-4'sd6))<<<((5'sd6)?(4'd1):(-3'sd3))))));
  localparam [3:0] p6 = (&{3{{2{(4'sd1)}}}});
  localparam [4:0] p7 = (~|{(-((5'sd7)?(3'd1):(4'd9))),{4{(4'sd7)}},((-3'sd1)?(4'd3):(-2'sd1))});
  localparam [5:0] p8 = (2'd2);
  localparam signed [3:0] p9 = ((((2'sd0)<<<(-4'sd3))*((-3'sd3)!==(-5'sd13)))>>>(^(~^(^(|(5'sd9))))));
  localparam signed [4:0] p10 = {3{({4{(2'd2)}}?{2{(3'sd0)}}:{1{(-3'sd0)}})}};
  localparam signed [5:0] p11 = (3'd4);
  localparam [3:0] p12 = (((5'd4)/(4'd9))?((2'sd0)?(3'd0):(5'sd7)):((-5'sd4)?(3'd1):(2'd3)));
  localparam [4:0] p13 = ((2'd3)!==(5'd21));
  localparam [5:0] p14 = ((((5'sd13)>=(5'd5))|((4'd3)<(4'd0)))<=(((-4'sd3)!=(5'd31))%(-3'sd1)));
  localparam signed [3:0] p15 = {((-5'sd0)^(5'd3)),((3'sd2)-(2'd2)),((4'd5)<<(5'sd14))};
  localparam signed [4:0] p16 = (2'd0);
  localparam signed [5:0] p17 = {4{{2{(4'sd2)}}}};

  assign y0 = (5'd24);
  assign y1 = (^(5'd2 * (p0-p2)));
  assign y2 = (~(|(~(|(&(+(~^(~|(&p7)))))))));
  assign y3 = (p10&p17);
  assign y4 = (~&({(~&b1),(p1&p7),(p17|b4)}+({{a2,b1}}<<(|{p17}))));
  assign y5 = (((^{{4{{2{(~p10)}}}}})));
  assign y6 = {{p15,p1,a3},{a0,p9,a4},(~{a0,a4,b0})};
  assign y7 = (5'd31);
  assign y8 = (^{4{((+p12)-(~|p14))}});
  assign y9 = ((((b4+p13)<<<{2{p3}})<(^(p16+p14)))<((~|(a2+a4))<={1{(b3-p17)}}));
  assign y10 = (4'd4);
  assign y11 = ({1{{p8,p11}}}>(2'd0));
  assign y12 = ((-2'sd1)?{1{(b3||a1)}}:((b4||a3)<<<(a5?a2:b2)));
  assign y13 = (+(5'd30));
  assign y14 = $signed((((|a2))?(b2?b3:p1):$unsigned({4{a0}})));
  assign y15 = (((~|{p1,p11,b2})));
  assign y16 = (b5===b4);
  assign y17 = ((-2'sd1)?(4'd6):(~&p13));
endmodule
