module expression_00496(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((!(3'd5))&(~&(-4'sd3)));
  localparam [4:0] p1 = (-((-(|(2'd0)))|(|((2'sd0)<(5'd8)))));
  localparam [5:0] p2 = ((4'd5)<<(5'd10));
  localparam signed [3:0] p3 = (((-4'sd3)?(2'd3):(-4'sd7))?((2'd3)?(5'd25):(-2'sd1)):((4'sd5)?(-5'sd11):(3'sd1)));
  localparam signed [4:0] p4 = ((4'd5)<<<({((2'sd1)?(-5'sd0):(4'sd7))}>((3'd0)<<(-3'sd0))));
  localparam signed [5:0] p5 = (((-4'sd4)^(5'sd2))?((2'd2)<<<(-4'sd3)):(5'd15));
  localparam [3:0] p6 = (~(!(-5'sd2)));
  localparam [4:0] p7 = (^((5'd27)>=(3'd1)));
  localparam [5:0] p8 = (4'd11);
  localparam signed [3:0] p9 = (((3'd7)>=(5'd24))!=((2'd1)-(5'sd8)));
  localparam signed [4:0] p10 = ((((-2'sd0)?(-4'sd2):(-2'sd1))&&(-(3'd7)))?(+((-2'sd1)!==(-3'sd3))):(-2'sd1));
  localparam signed [5:0] p11 = (((3'd0)-(-4'sd6))<<((5'd3)?(-5'sd1):(5'd18)));
  localparam [3:0] p12 = (4'd10);
  localparam [4:0] p13 = (^(~|((~|(-3'sd0))?(~(-3'sd0)):(~|(-4'sd4)))));
  localparam [5:0] p14 = ((5'd1)^~(3'd7));
  localparam signed [3:0] p15 = ((2'sd0)?(-3'sd0):(2'd0));
  localparam signed [4:0] p16 = {((5'sd10)>>(2'd3)),{(4'd12)},{(2'sd0),(2'd3)}};
  localparam signed [5:0] p17 = ((-2'sd1)?((-5'sd13)==(4'd8)):(+((5'd3)^(-2'sd0))));

  assign y0 = (4'd7);
  assign y1 = ({4{p0}}<={4{b2}});
  assign y2 = (2'sd1);
  assign y3 = ($signed(((~&b5)!==(b2>=a2)))>>((-2'sd0)?(!p9):(|a4)));
  assign y4 = (^(+{2{{1{{3{(~&{3{p13}})}}}}}}));
  assign y5 = ((a0?p4:b1)>>>($signed((~&p0))));
  assign y6 = {((b0+b4)===(2'd2)),{{b0,a3},{a3},(a1?p5:b0)},((5'd9))};
  assign y7 = (((-(b4<p17))!=(-2'sd1))>>((-(b3===a2))>{3{a0}}));
  assign y8 = $unsigned({$signed(p3),(b5<<p2),{3{a0}}});
  assign y9 = ({(a3===a5),(2'd1),(p1?a3:a4)}||(!((p7<p4)?{1{p0}}:(~|p1))));
  assign y10 = (3'sd3);
  assign y11 = (((a0?p10:a2)?(a2+a2):{a1})-{(a2==a5),(a1?a0:b3)});
  assign y12 = $unsigned((4'd1));
  assign y13 = ((a2?p2:a4));
  assign y14 = (((p5?p0:p6)?(p12?p2:b5):(p13?p4:p4)));
  assign y15 = (+(-(((5'd22)==(a3?p2:a2))|(-3'sd2))));
  assign y16 = ({2{(p15>=a1)}}<<({3{p3}}?{2{p0}}:(-p0)));
  assign y17 = (5'd2 * (b0?p2:p2));
endmodule
