module expression_00566(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{2{(5'd4)}}}};
  localparam [4:0] p1 = ((+(-3'sd1))%(2'd2));
  localparam [5:0] p2 = ((5'd4)&(3'sd3));
  localparam signed [3:0] p3 = ((3'sd3)&(-4'sd0));
  localparam signed [4:0] p4 = ({(3'd0)}?{(2'sd0)}:{(3'sd0)});
  localparam signed [5:0] p5 = {2{{2{(2'sd0)}}}};
  localparam [3:0] p6 = ((((5'd2)<(-5'sd0))&((4'sd4)!==(-4'sd4)))?((~&(3'sd0))?(2'd2):(~|(3'd5))):((-(3'sd0))*(^(3'd5))));
  localparam [4:0] p7 = {2{{4{{2{(-5'sd10)}}}}}};
  localparam [5:0] p8 = (((^((4'sd6)>>(4'd12)))<((-4'sd2)<(4'd4)))>>(4'sd4));
  localparam signed [3:0] p9 = (-5'sd8);
  localparam signed [4:0] p10 = (-5'sd1);
  localparam signed [5:0] p11 = (|(^(|((&(4'sd1))==((5'sd14)|(5'd29))))));
  localparam [3:0] p12 = ((((5'd22)?(5'd21):(2'd2))?((5'sd11)-(2'sd1)):((3'd0)?(5'd27):(4'd9)))>=({(4'd11)}>>>((4'd3)>>>(-4'sd6))));
  localparam [4:0] p13 = {3{(&((5'sd13)===(5'd12)))}};
  localparam [5:0] p14 = ((~|((3'd5)^~(3'sd2)))>=((3'd0)!==(2'd2)));
  localparam signed [3:0] p15 = ({2{(5'd11)}}?((3'd6)<(4'd3)):(!{4{(-5'sd0)}}));
  localparam signed [4:0] p16 = ({(((4'sd7)?(3'd1):(4'sd3))?{1{(2'sd0)}}:{(4'sd5)})}|({4{(5'd31)}}!==((-5'sd2)?(2'd0):(5'sd0))));
  localparam signed [5:0] p17 = (+(2'sd1));

  assign y0 = (&(^(^(-3'sd1))));
  assign y1 = ((a4?a5:p12)*(a5<<<p4));
  assign y2 = ({(p5?p0:p1),(a1?p7:p7),{(a1===a2)}}>>((p15?p13:p9)?{a2,p6,p5}:(6'd2 * b0)));
  assign y3 = ((3'sd2)?{1{(3'd0)}}:{(2'd2),{a4,b3,b1},(b5?p9:p15)});
  assign y4 = (-(~|((5'sd14)<<((|(p6>>p9))?(4'sd6):(p17<=p3)))));
  assign y5 = (~|(((b5?b3:b3)>(a4===b0))<<<$unsigned((a1?a2:b4))));
  assign y6 = ((~^p7)&&{b4,p15,p2});
  assign y7 = (b2<<<p11);
  assign y8 = (({4{p14}}<<(p12?b1:p2))&&({3{p16}}?(p1?p14:b0):(p13?p10:p8)));
  assign y9 = {{(p2?p15:p14),{(p9!=p17),(b2?b1:b1)}}};
  assign y10 = {{((a1^~a3)>{a1,b4}),({(a2>=a5)}!=(a1^a4))}};
  assign y11 = $unsigned((~$signed(((((4'd8)%p8)<<((b4<<<p14)))<<(((~^a0)<(a1===a1))||(~(-$unsigned(a5))))))));
  assign y12 = (({4{p13}})>(~|(~(3'sd0))));
  assign y13 = (~(5'd16));
  assign y14 = (p10==p9);
  assign y15 = {{{{p9},{p8}}},{{p0},{p2}},{{p0},{a5}}};
  assign y16 = $signed((((p13?p1:p6)/p1)?((p8&&p17)*(b3?p14:p8)):((p8-p8)<=(p17?p1:p4))));
  assign y17 = (b3?b3:p13);
endmodule
