module expression_00526(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd2)-(3'sd1))/(2'd1));
  localparam [4:0] p1 = (|((((5'd23)^~(3'd3))|((-4'sd0)!=(5'sd10)))>=(-((!(5'sd9))==(4'd10)))));
  localparam [5:0] p2 = (-{3{(-(!((2'd2)!=(2'd1))))}});
  localparam signed [3:0] p3 = (&(4'd4));
  localparam signed [4:0] p4 = (((5'sd4)^~(2'sd1))<((3'd7)&&(5'd5)));
  localparam signed [5:0] p5 = {(3'sd3),(~&(2'd3))};
  localparam [3:0] p6 = {{(&(4'd3)),((~&(4'd0))?((-4'sd1)?(3'sd0):(-5'sd12)):(-2'sd1))}};
  localparam [4:0] p7 = ((4'd3)|(-3'sd0));
  localparam [5:0] p8 = ((+(4'd2 * ((4'd11)<<(2'd3))))<=((~^((3'sd3)^~(3'd5)))&&(-(~^(~|(-4'sd3))))));
  localparam signed [3:0] p9 = ((3'd4)?{1{((-3'sd0)?(-2'sd0):(4'sd3))}}:(|((3'd3)?(5'sd15):(-2'sd0))));
  localparam signed [4:0] p10 = {{(4'd2 * ((3'd4)+(4'd14)))},(-3'sd1)};
  localparam signed [5:0] p11 = (~(5'd11));
  localparam [3:0] p12 = ((3'sd2)&&(3'd6));
  localparam [4:0] p13 = ((4'd9)>=(((4'sd4)==(2'd1))<<<((3'sd2)>=(-2'sd0))));
  localparam [5:0] p14 = {3{(~((5'd17)?(-3'sd0):(-2'sd0)))}};
  localparam signed [3:0] p15 = (&(3'sd1));
  localparam signed [4:0] p16 = {4{((4'd10)|(5'd1))}};
  localparam signed [5:0] p17 = (((5'd3)?(4'd11):(2'd2))?((3'sd2)!==(2'd1)):((2'd1)?(5'sd2):(2'd1)));

  assign y0 = ((5'd26)<<<(2'd2));
  assign y1 = (3'd6);
  assign y2 = {4{(p3?p4:p14)}};
  assign y3 = (({a1}<(b1?p11:b2))?({b3,b1}^~{a4}):{(p2<=a4),{p0,a2},(b4||p14)});
  assign y4 = ((((p12!=a5))-(+(4'sd7)))!=$signed((~&(|((b0?b0:a1)==(|b0))))));
  assign y5 = (!$signed(((2'sd0)?$unsigned((~(4'd0))):$signed($signed((-3'sd2))))));
  assign y6 = {1{(~^((~&(~^(p2?b3:b3)))>>>({2{p5}}?(b3?b1:p3):(!a3))))}};
  assign y7 = (~&((~&(~&(+(&{(!b0),{p2,p10,a1}}))))<{(~{b4,p7}),(!(+(6'd2 * p12)))}));
  assign y8 = (+$signed({({a5,p5}),(p13||b5)}));
  assign y9 = (-5'sd10);
  assign y10 = (2'sd1);
  assign y11 = {(^{2{{(+(&{p0,p14,a5}))}}})};
  assign y12 = {{4{p2}},{b4,a0,p4},((a5?b0:b2)>(b4>p17))};
  assign y13 = ({3{p3}}>=(!(b0===a4)));
  assign y14 = ((|((+(b0<b5))<(~(b2&a1))))&((!(a4!=b2))<=(b3*b3)));
  assign y15 = (((a1&&b0)||(p15^p14))>((p17-a5)-(a4>=b4)));
  assign y16 = {3{{2{p15}}}};
  assign y17 = {2{((~{3{p3}})&&(2'd1))}};
endmodule
