module expression_00730(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-2'sd1);
  localparam [4:0] p1 = ((((4'sd3)?(5'd15):(-5'sd13))?((5'd30)?(3'sd3):(5'd7)):{(3'd0),(-5'sd10)})?({(3'd6),(2'd2)}?{(-4'sd4),(-5'sd9),(-2'sd1)}:{(-2'sd0),(-5'sd5),(2'd3)}):(((3'd1)>>(-4'sd2))^{(3'd1)}));
  localparam [5:0] p2 = (5'd25);
  localparam signed [3:0] p3 = (~^(^(~^{(-({{((-5'sd1)>>(2'd0))}}==((5'd2 * (3'd2))===(4'd7))))})));
  localparam signed [4:0] p4 = (!{4{(!(3'd4))}});
  localparam signed [5:0] p5 = ({(-(((3'd0)===(-5'sd11))^~(!{(3'sd3)})))}>=((((5'd14)!=(4'sd2))^((4'd8)-(-5'sd14)))===(+((-3'sd3)?(-4'sd7):(3'd3)))));
  localparam [3:0] p6 = (!{(&(4'sd7))});
  localparam [4:0] p7 = ((~^{((3'sd2)?(-5'sd5):(-2'sd0)),(~(2'd0))})>={4{(4'd9)}});
  localparam [5:0] p8 = (((~^(-4'sd1))^~((-2'sd1)?(3'd7):(-2'sd1)))<=(((5'sd8)?(3'd7):(-4'sd4))?((4'd13)&(4'd13)):((4'd12)&(-2'sd0))));
  localparam signed [3:0] p9 = (-((-5'sd8)?(2'd2):(2'sd0)));
  localparam signed [4:0] p10 = (+((|((-4'sd6)%(5'd4)))|((~&(4'sd0))<<(-(4'sd6)))));
  localparam signed [5:0] p11 = (((^{(4'd8)})>>((5'd9)&(2'sd0)))=={(4'd7),(-4'sd3)});
  localparam [3:0] p12 = (~&{(&(~|({2{(-4'sd6)}}>>>{(5'd7),(3'sd1)})))});
  localparam [4:0] p13 = {(!{(5'd8),(3'sd0)}),(+(|(-4'sd5)))};
  localparam [5:0] p14 = ((((^(2'd1))!=((3'sd3)>(3'sd1)))>{4{(2'd1)}})==(-{4{(6'd2 * (5'd7))}}));
  localparam signed [3:0] p15 = {3{(+{4{(-5'sd0)}})}};
  localparam signed [4:0] p16 = {3{(4'd7)}};
  localparam signed [5:0] p17 = (-(4'sd0));

  assign y0 = (({1{((p7==b4)>>(a4===b3))}}&{(4'd7)})>{(p16==b2),(~^{p9,p11,p1}),{3{b4}}});
  assign y1 = ((p2%a2)!=(b1!==a2));
  assign y2 = ((~(4'd2))/a2);
  assign y3 = ((a0===b4)>(b5%b3));
  assign y4 = (~^(a1^b1));
  assign y5 = (!b1);
  assign y6 = {((~^(&b1))?(b5?b4:p9):(!(p14?p16:p12))),{({a2,p15}?(b2?p6:p15):{(-b4)})}};
  assign y7 = (+(2'd2));
  assign y8 = (~((+(p12?p6:a4))?(a1?p11:a0):(a0?p2:a4)));
  assign y9 = {2{({3{p3}}<<<({4{p4}}))}};
  assign y10 = ((p16^p15)<=(p4-p5));
  assign y11 = (&(~a0));
  assign y12 = (((4'd2 * p2)>=(a2*a4))^((p2^p5)!=(a0|p9)));
  assign y13 = $unsigned($signed({p16,p5,a2}));
  assign y14 = ((&(&(5'sd3)))?((+((3'd2)?(b5):(2'd0)))):((4'd11)?(b4):(2'd1)));
  assign y15 = (p5>p5);
  assign y16 = ((a3?a1:a0)?((a0<b3)>=(5'd2 * a1)):((4'd2 * a2)+(a0?b0:a5)));
  assign y17 = {1{(5'd2 * (-(p2&p8)))}};
endmodule
