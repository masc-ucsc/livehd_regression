module expression_00375(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((6'd2 * ((3'd2)>>>(5'd4)))!=(((5'd22)+(2'd1))^~((-4'sd4)^(3'd6))));
  localparam [4:0] p1 = (-((2'd1)?(-4'sd4):(2'd1)));
  localparam [5:0] p2 = {((5'd2 * (~^(~&(4'd10))))<(((4'd13)+(5'd2))>((-3'sd3)>>(4'd11))))};
  localparam signed [3:0] p3 = ((((~&(4'd4))^~(&(2'sd0)))==(~&((-5'sd4)>>(4'd1))))>(((+(-3'sd3))<=(|(2'd3)))==(^(~^(-(2'd0))))));
  localparam signed [4:0] p4 = ((((4'd2)<<<(4'd4))|((3'sd1)<<<(5'd21)))>>>(((3'd6)||(3'sd0))<((2'sd1)*(-2'sd1))));
  localparam signed [5:0] p5 = (((2'd3)==(5'd6))?((4'd3)>(4'd6)):((2'd1)^(-4'sd6)));
  localparam [3:0] p6 = (({3{(5'd28)}}&&((3'd3)|(4'd15)))<(~^(~&{((5'd12)!==(3'd2)),{(3'd4)},((-2'sd0)>=(2'sd0))})));
  localparam [4:0] p7 = {3{{3{(2'd1)}}}};
  localparam [5:0] p8 = (({2{(3'd3)}}||{(5'd24),(-5'sd5)})&&{((2'd3)>=(4'd3))});
  localparam signed [3:0] p9 = ({4{(-2'sd1)}}>>>(-5'sd0));
  localparam signed [4:0] p10 = ((~|((-3'sd3)?(2'sd1):(5'sd14)))?((5'd11)?(3'd1):(3'd5)):(~&(~|(3'd5))));
  localparam signed [5:0] p11 = (((4'd0)&&(-5'sd15))&&(&((2'sd1)||(5'sd9))));
  localparam [3:0] p12 = {(-(&{{(3'sd1),(3'd5),(2'd3)},(-(3'd0)),((-5'sd10)?(-5'sd8):(2'd3))})),(-(!(^(&((5'd23)!=(-5'sd9))))))};
  localparam [4:0] p13 = {({(-3'sd1),(5'sd13),(-2'sd1)}>={(2'd0)}),({(4'd1),(-5'sd1),(4'd5)}<{(4'd13)}),{({(2'sd1)}<{(-5'sd3),(5'sd14),(-3'sd3)})}};
  localparam [5:0] p14 = (((6'd2 * (3'd7))+((4'd8)<<<(-3'sd1)))<<{((3'd7)>(3'd4)),((5'd18)>=(2'd0))});
  localparam signed [3:0] p15 = ((5'd3)^~(-2'sd0));
  localparam signed [4:0] p16 = ((!((~|(-3'sd0))&&(-(2'd3))))||((~&(-(2'd3)))<<((4'd0)*(-2'sd0))));
  localparam signed [5:0] p17 = (-4'sd1);

  assign y0 = (|a3);
  assign y1 = (!(~(~&{2{((~p10)>>>(a0>>b3))}})));
  assign y2 = ({1{{4{p8}}}}?({1{a5}}>>{b2,p10}):({4{p11}}<=$signed(p15)));
  assign y3 = ((b0||a5)<={1{(~^a0)}});
  assign y4 = ($unsigned(($signed(p6)?$unsigned(b0):(a3)))>>>(((a0>b5)^(p8?b5:b1))||(a5?a3:p13)));
  assign y5 = ((|(^{$signed((!((b5)<{b2,a2})))}))!=={(5'd2 * {3{b2}}),{{4{a2}},{a0,b3},{2{a4}}}});
  assign y6 = (2'd1);
  assign y7 = {(~|(4'd2 * {(p13>p2)}))};
  assign y8 = (~{(2'd1),(-{p2,p4}),(5'sd10)});
  assign y9 = {1{{3{({2{b1}}>{1{p8}})}}}};
  assign y10 = {((b3^~a4)^(b3!=b3)),{(b0?b1:b2),{p9,p8,p2}},((b0?b2:p16)>{p10,p9})};
  assign y11 = (-4'sd5);
  assign y12 = (((p8==a3))>((p13+a1)));
  assign y13 = (!{(p3&b5),{p4,a5},(a5<<a5)});
  assign y14 = {4{a3}};
  assign y15 = (({(&{4{b0}}),(4'sd1)})!=(!(^((3'sd1)&(5'd29)))));
  assign y16 = {4{((a5<=p5)>$unsigned(a0))}};
  assign y17 = (^$signed((~|(~$signed($signed(($unsigned({(!p3),$signed(p9)})>=(~^{$unsigned(b2),(|p9),$signed(p11)}))))))));
endmodule
