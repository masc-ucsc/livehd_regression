module expression_00458(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(+(5'sd7)),(~&(5'sd12))};
  localparam [4:0] p1 = (~&(((-4'sd4)?(-4'sd7):(4'd8))?((2'd3)?(4'd15):(2'd1)):(2'd2)));
  localparam [5:0] p2 = (5'd9);
  localparam signed [3:0] p3 = ((-2'sd1)<(5'd24));
  localparam signed [4:0] p4 = {(~&(!(~(4'd10)))),({(3'd4),(4'sd1),(2'd3)}>{(4'd9),(5'sd14)}),(!(^((3'd7)===(4'sd0))))};
  localparam signed [5:0] p5 = ((-4'sd2)?{((-3'sd1)?(5'd18):(2'd2))}:{4{(-4'sd4)}});
  localparam [3:0] p6 = (((5'sd13)?(4'sd1):(3'd4))?{1{(-4'sd0)}}:(-4'sd4));
  localparam [4:0] p7 = ((((4'sd1)?(-3'sd1):(4'd8))+((-4'sd0)?(2'sd0):(-2'sd0)))?(((-4'sd5)||(4'sd4))*((5'd4)?(3'd3):(3'sd2))):(((-5'sd1)>=(2'sd0))+((5'sd0)&(5'd11))));
  localparam [5:0] p8 = (+(~|((^((4'd8)||(2'd3)))+(~{2{(-2'sd1)}}))));
  localparam signed [3:0] p9 = (4'd2 * (2'd2));
  localparam signed [4:0] p10 = {(5'sd11),{{3{(-4'sd7)}}},((2'sd0)+{(3'd3),(2'd3),(2'sd1)})};
  localparam signed [5:0] p11 = ((((3'd0)?(2'd1):(-5'sd4))?(|(2'd1)):((-4'sd3)?(-3'sd1):(4'd8)))?(((3'sd0)?(2'd2):(-3'sd3))>=(^(-5'sd2))):((+(3'sd1))?((4'sd7)<<(-2'sd0)):(~|(-5'sd14))));
  localparam [3:0] p12 = (((4'd9)==((-3'sd0)+(4'd5)))>>>((((5'd26)==(4'd12))<<<((4'd6)>=(5'd16)))>>>(6'd2 * ((3'd0)%(4'd13)))));
  localparam [4:0] p13 = {{(5'd27),(3'sd1),(3'd0)}};
  localparam [5:0] p14 = (2'd1);
  localparam signed [3:0] p15 = {{(2'sd1),(3'sd1),(2'sd1)},{(-2'sd1),(4'd13),(2'sd0)},{(3'd4),(-2'sd1),(-3'sd3)}};
  localparam signed [4:0] p16 = ({(3'sd3),(3'sd0),(5'd6)}+{4{(-5'sd5)}});
  localparam signed [5:0] p17 = (3'd7);

  assign y0 = ({1{(({3{a3}})<<{1{(3'd6)}})}}&&(2'sd1));
  assign y1 = ((~^((+p17)?(-p10):(p7)))>>((p16?a5:p17)>>(!(p3?p6:b4))));
  assign y2 = {4{({4{p9}}&(p11>=p14))}};
  assign y3 = (4'd0);
  assign y4 = {2{(4'd8)}};
  assign y5 = (((5'd15)&(b1?a2:p14))-((b0<=a0)?(a4&&a2):(a5&b5)));
  assign y6 = (~&(~(~{a4,a2,p1})));
  assign y7 = (4'd8);
  assign y8 = $signed({2{b4}});
  assign y9 = (!(p17-p16));
  assign y10 = (&((b3>>p10)<=(^(^b0))));
  assign y11 = (((~|(+p8))>={p8,p7})>>{(~(a3===b2)),(+(a0^b4))});
  assign y12 = ((!((~^(~(a0?b2:b3)))+(+(a5==b4))))>=(~(~&(^(+((b3!=a5)*(6'd2 * b2)))))));
  assign y13 = {{3{{2{{2{p14}}}}}}};
  assign y14 = (&(((a5!==b4)||{2{p9}})>(-{1{(p8>>>p13)}})));
  assign y15 = {4{(&(3'sd3))}};
  assign y16 = ({(-4'sd6),(-5'sd10),{(p6>>>a2)}}&&((5'd2 * (5'd28))&&((5'd1)>=(b1&a3))));
  assign y17 = ((!(^(p3?a4:b1)))<<<$signed((a0<<a1)));
endmodule
