module expression_00560(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-((-5'sd15)^~{{1{(4'd4)}},(5'sd15),(2'd0)}));
  localparam [4:0] p1 = (5'd13);
  localparam [5:0] p2 = {1{((-{3{(4'd7)}})<=((3'sd3)==(4'sd1)))}};
  localparam signed [3:0] p3 = {1{{4{((3'd6)!=(5'd19))}}}};
  localparam signed [4:0] p4 = {3{{3{(3'd5)}}}};
  localparam signed [5:0] p5 = (!(+{3{(5'd2 * (2'd0))}}));
  localparam [3:0] p6 = ({4{(2'd2)}}?(-5'sd8):(((-5'sd6)?(5'd25):(2'sd1))&((3'd1)?(4'd12):(5'sd13))));
  localparam [4:0] p7 = (((5'd31)?(2'd1):(3'd0))?(((5'd18)>>(3'd5))&(3'd0)):{4{(2'd1)}});
  localparam [5:0] p8 = ((((-4'sd2)>(-3'sd2))!=(4'sd5))>>>{(2'd1),(-3'sd2),(2'sd1)});
  localparam signed [3:0] p9 = (^(~((2'd2)<(-2'sd1))));
  localparam signed [4:0] p10 = ((((4'd1)&&(2'd1))+((2'd2)==(2'sd0)))?({2{(5'sd3)}}^(|(4'd13))):((4'd2 * (2'd3))&((-3'sd2)?(4'd12):(3'd3))));
  localparam signed [5:0] p11 = ((^(5'sd11))|{2{(-2'sd1)}});
  localparam [3:0] p12 = (((4'sd7)?(5'sd14):(4'd10))=={3{(2'd1)}});
  localparam [4:0] p13 = {{({(&(-2'sd1)),((5'sd4)||(2'sd0)),{(-2'sd1),(3'd2),(2'd2)}}!=={(-((4'd4)?(3'd5):(3'd4))),((4'd9)^~(3'd7))})}};
  localparam [5:0] p14 = (+((~^(+(((3'd5)!==(3'd7))!=((3'sd0)-(2'sd0)))))>>((-((2'd3)%(-2'sd1)))^((2'd2)*(5'd30)))));
  localparam signed [3:0] p15 = {((4'sd6)-(3'sd0)),((4'd2)-(3'd5))};
  localparam signed [4:0] p16 = ({2{(2'd1)}}?(5'd28):{3{(-2'sd1)}});
  localparam signed [5:0] p17 = ((~&(&(-5'sd2)))+(~|(&(4'd10))));

  assign y0 = {((p15^~p2)<<{p1}),{((p4&p10)^~(p1?p5:p3))}};
  assign y1 = (&{((^(|p12))^~(b3>=b3)),{(b3==a3),{p17},{p3,b5}}});
  assign y2 = (((~|p3)?(p13<<p4):(-p10))<<<({2{p7}}&$unsigned(a0)));
  assign y3 = ((p15?b1:p7)^~((p6<=p8)&{p17}));
  assign y4 = (~&{(~|(!(~({b3,a5}^{a5})))),((b3===b0)?(!a5):(2'sd1))});
  assign y5 = $signed((((b3?b2:a0)+((a2&&a5)^~(a0<a4)))&((b0?p11:p3)&&{b0,b2,p16})));
  assign y6 = (^((~&((~^p14)?(^p6):(^p13)))&&((|(&p6))/p15)));
  assign y7 = {4{{2{{3{b3}}}}}};
  assign y8 = ((($unsigned(($signed(a5)?(a3!==b1):(b1===a1)))))<=(((b2>>>b1)+(b3?b2:p14))<=(b3?p16:b4)));
  assign y9 = ((p17?p16:p16)?(5'sd14):(+p17));
  assign y10 = {3{(a1<<p12)}};
  assign y11 = {4{{3{p5}}}};
  assign y12 = (~|(&(&(-(~&((~^(+(~((a4|a0)&(~a1)))))>=((p15>>b3)*((+b4)))))))));
  assign y13 = (+p16);
  assign y14 = ((b1*b4)+(b5>b3));
  assign y15 = ({3{{3{{1{p0}}}}}});
  assign y16 = $unsigned(((p17&p11)^~((b5&p4))));
  assign y17 = {{{b1,p8}},{{b4,a1,b5},{b4}}};
endmodule
