module expression_00633(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((((-2'sd1)%(2'sd0))&&((5'd14)-(2'sd1)))>((~&(5'sd11))>=(-(4'sd7))))||(((!(4'sd5))>>((-2'sd0)<<(3'd5)))-((|(2'sd0))+((2'sd1)|(4'd15)))));
  localparam [4:0] p1 = (^(~&(5'd28)));
  localparam [5:0] p2 = (~^(-5'sd5));
  localparam signed [3:0] p3 = ((3'd7)?(3'sd0):(2'sd1));
  localparam signed [4:0] p4 = (((4'd5)?(2'd1):((-5'sd14)&(4'sd6)))<<{3{((-4'sd3)||(4'd3))}});
  localparam signed [5:0] p5 = (({2{(-3'sd1)}}<<<{(-5'sd13),(2'd3),(4'd4)})<=({4{(3'd4)}}!={3{(-4'sd2)}}));
  localparam [3:0] p6 = {2{{1{{2{(-4'sd6)}}}}}};
  localparam [4:0] p7 = {(~^{(3'd2),(4'd9),(4'sd7)}),(~^{2{(3'sd0)}}),(~^(&(-5'sd4)))};
  localparam [5:0] p8 = ((5'd14)?(3'd0):(5'd20));
  localparam signed [3:0] p9 = {4{(4'd5)}};
  localparam signed [4:0] p10 = (^(((^(3'd2))?(~^(5'd27)):((3'sd3)&&(3'd6)))?((~|(2'd0))?(6'd2 * (4'd13)):((3'd3)?(-4'sd2):(4'sd1))):(~&(~^((5'd13)!=(4'd3))))));
  localparam signed [5:0] p11 = (&((3'd6)>>(2'sd0)));
  localparam [3:0] p12 = (((-5'sd1)?(5'sd9):(5'sd4))==((4'sd6)?(4'd8):(2'd2)));
  localparam [4:0] p13 = ((!({((-5'sd7)>>>(-5'sd6))}&{2{(5'd11)}}))+(!({1{(+(5'sd14))}}&&((-5'sd3)!=(4'd7)))));
  localparam [5:0] p14 = (((4'd5)?(-3'sd1):(5'd10))<<<{((5'd2)>>>(3'd4))});
  localparam signed [3:0] p15 = ((5'd19)?(|(-3'sd0)):(5'd15));
  localparam signed [4:0] p16 = (((3'd2)>(2'd0))>>(5'd8));
  localparam signed [5:0] p17 = {4{{1{(3'sd0)}}}};

  assign y0 = {4{((p4?p1:a4)?(p14?p1:b0):(p10|p3))}};
  assign y1 = (-{(a5<=p7),(p10<=a5),(p6>>>p6)});
  assign y2 = (5'd6);
  assign y3 = ({3{(b3<<p8)}}>>(|(!((p13||p1)))));
  assign y4 = {3{((^a1))}};
  assign y5 = {((p3?p7:p17)||(|{p12,p17}))};
  assign y6 = (|(((b5?b3:a4)?(-(a0-b0)):(a0!==b1))|(5'd25)));
  assign y7 = (+(((!b2)?(~&a3):(a2?b4:b5))>=(((p3^a2)/a4))));
  assign y8 = {$signed(b0),$signed(b2),$unsigned(b0)};
  assign y9 = ({(5'd2 * (^p0)),(|(p12<<<p6))}<=((~|$unsigned($signed(b0)))!=={2{{2{a5}}}}));
  assign y10 = {3{(b2<=a1)}};
  assign y11 = ((^p15)?$unsigned(p15):(&p5));
  assign y12 = {1{(((a5!=p1)<<(p6>p7))>((p16<<p4)>=(4'd2 * p6)))}};
  assign y13 = ((a4?b0:p11)?(p15?p12:p8):{(-a2)});
  assign y14 = (~^(!(|((((-4'sd6)<<(|b1)))^(~(4'sd6))))));
  assign y15 = (2'd3);
  assign y16 = (+(5'sd4));
  assign y17 = (((~(p3>a1)))==$signed((~^$unsigned({p11,p8}))));
endmodule
