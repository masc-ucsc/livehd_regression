module expression_00969(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd12)?(5'sd15):(2'd0))?(-4'sd5):(2'sd1))||(4'd2 * ((3'd4)/(4'd5))));
  localparam [4:0] p1 = (-{3{{1{(3'd6)}}}});
  localparam [5:0] p2 = {{{(2'd0)},{(5'd5)}},({(3'sd3),(-4'sd3),(-4'sd4)}<{(3'sd1),(4'sd2)})};
  localparam signed [3:0] p3 = ((&((2'sd1)>=(3'd2)))<(2'd3));
  localparam signed [4:0] p4 = ((2'd1)>>{{(4'd6),(3'd1)}});
  localparam signed [5:0] p5 = {4{((-2'sd0)>>>(-3'sd3))}};
  localparam [3:0] p6 = ((((-3'sd3)^(2'd3))>=((4'sd3)===(5'sd15)))+({2{(-4'sd6)}}===((3'sd3)&(2'd1))));
  localparam [4:0] p7 = (((~&(2'd2))<((-5'sd6)<<(-5'sd5)))!==(((-4'sd4)<(2'd1))<<<((5'sd5)?(-4'sd7):(5'd9))));
  localparam [5:0] p8 = (5'd10);
  localparam signed [3:0] p9 = ({(2'sd1),(3'sd3),(4'd6)}?(-(6'd2 * (2'd2))):{(-3'sd1),(5'd7),(2'd0)});
  localparam signed [4:0] p10 = ((2'd0)?((3'd7)?(4'sd7):(3'd3)):(((5'sd1)?(5'sd14):(4'd1))<<((-2'sd0)?(3'd3):(-4'sd3))));
  localparam signed [5:0] p11 = (~|(4'd10));
  localparam [3:0] p12 = (!(|{4{(-5'sd14)}}));
  localparam [4:0] p13 = ((4'd10)?(2'd2):(4'd12));
  localparam [5:0] p14 = {{{(3'd4)},{(-3'sd0),(-4'sd5)}},{(2'sd0),(4'd6),(4'd11)}};
  localparam signed [3:0] p15 = {((|(-2'sd1))?((5'sd15)>(4'd4)):(&(-5'sd11))),(((-2'sd1)?(-4'sd2):(3'd6))-((-2'sd0)>>>(2'sd1))),(-((2'sd0)?(4'd0):(5'sd10)))};
  localparam signed [4:0] p16 = {4{(!((2'sd1)<=(4'd13)))}};
  localparam signed [5:0] p17 = ((((5'sd10)|(-2'sd1))>>((3'sd2)?(4'd9):(5'd1)))>>>{3{((3'sd3)^~(2'd3))}});

  assign y0 = ((((b4-a3)<<<(b0?b5:a0))-((-b3)<=(a1?b5:a1)))===((a1?b5:a4)?(b4?b3:b1):(b0||b0)));
  assign y1 = (4'd14);
  assign y2 = ((-5'sd1)&(^((^p15)?(5'd20):{4{p5}})));
  assign y3 = ((p8*p8)/p0);
  assign y4 = (-(((a4?a1:a0)?$unsigned(b2):(a0?a1:p17))<<<((&b5)?(b4<<<p16):(a4-a2))));
  assign y5 = {(4'd7),(-(3'd2))};
  assign y6 = ((p13?p7:p8)?$signed(p13):(a3<<a3));
  assign y7 = (({1{(2'd1)}}|(a4&&b0))&(5'd4));
  assign y8 = $signed({2{{4{{3{a2}}}}}});
  assign y9 = ((p13)<<(p15+p8));
  assign y10 = ({1{(|((b2?p4:a0)))}}?({2{p10}}?(a3!=p2):(b0&&p15)):((-b5)?(a4?b3:p12):(b0?p13:p6)));
  assign y11 = ((+{(p8>>>b3),(5'd2 * p0)})?(-{(+(a0^p0)),(-(-a1))}):((p1?b1:a0)?{a0,b3}:{p9}));
  assign y12 = (&(((!p5)?(b2):(-p2))<<<$signed((6'd2 * (-(^a2))))));
  assign y13 = {3{p2}};
  assign y14 = ((b3?b4:a4)^~{1{(5'd2 * b1)}});
  assign y15 = {((6'd2 * a0)^~(b0?a4:b1)),((b2>=b4)?(-5'sd11):{a1})};
  assign y16 = (2'd1);
  assign y17 = (($signed((-5'sd4))===(5'd28))<<((4'd3)));
endmodule
