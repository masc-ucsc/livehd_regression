module expression_00525(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(&(-((!((5'd7)-(5'sd15)))<=((|(5'd15))==((5'sd9)^~(3'd2)))))));
  localparam [4:0] p1 = (-5'sd4);
  localparam [5:0] p2 = ((((4'sd1)&(-4'sd4))<=((3'd6)/(4'd4)))+(((4'sd4)||(-4'sd4))==((-2'sd0)||(3'd2))));
  localparam signed [3:0] p3 = {{(2'sd0),(-2'sd0)},((3'd5)?(5'd24):(5'd13))};
  localparam signed [4:0] p4 = {{((((4'd8)==(3'd7))==((2'd1)>>(5'd31)))==={{(4'd7)},((3'd7)>=(3'd0)),((4'sd1)>(-2'sd0))})}};
  localparam signed [5:0] p5 = (((5'sd14)?(-3'sd0):(2'd2))?((4'd15)?(-2'sd1):(2'd1)):((5'sd10)?(2'd1):(5'd8)));
  localparam [3:0] p6 = (+(-2'sd0));
  localparam [4:0] p7 = ((-2'sd1)?(5'd28):((5'd7)?(3'd6):(-4'sd7)));
  localparam [5:0] p8 = (~|(~|(3'd1)));
  localparam signed [3:0] p9 = {1{(-2'sd0)}};
  localparam signed [4:0] p10 = {1{(-3'sd1)}};
  localparam signed [5:0] p11 = ((2'sd1)?(5'd22):(-3'sd1));
  localparam [3:0] p12 = (((-4'sd1)?(5'sd8):(4'sd1))&&((3'd2)?(2'd2):(-5'sd13)));
  localparam [4:0] p13 = (~&(+(|{2{{3{(3'd3)}}}})));
  localparam [5:0] p14 = ((((3'd5)+(5'sd15))>>(!(-5'sd6)))?(((4'd7)<<(3'd3))?((5'd24)?(3'd1):(4'd2)):((4'd2)?(4'd7):(2'd1))):(((4'd2)?(-2'sd1):(4'sd6))<=((5'd8)>>>(4'd8))));
  localparam signed [3:0] p15 = ({3{{1{((3'sd1)>>>(-5'sd3))}}}}!=({2{{1{(-5'sd12)}}}}>{3{(3'sd0)}}));
  localparam signed [4:0] p16 = {1{(((4'd5)>=(-5'sd7))-(!(|(5'd12))))}};
  localparam signed [5:0] p17 = {{2{{4{(-4'sd4)}}}},{3{{(2'sd1)}}},{3{{1{(-2'sd0)}}}}};

  assign y0 = {(b5?b1:p0),((p9^~b5)<=(4'd8)),(a2?b5:a0)};
  assign y1 = ($signed(a5)?{a4}:(b2));
  assign y2 = ((&((~(6'd2 * b1))>=(~|(5'd8))))<((4'd5)>=(-(~(b5*b1)))));
  assign y3 = (b5||a2);
  assign y4 = (b3?p5:p3);
  assign y5 = {3{{((&b5)||(b4^~b5))}}};
  assign y6 = (p3-p5);
  assign y7 = ((5'd2 * (a1!==a0))-$signed(((a2))));
  assign y8 = (((p5^~p1)|(p12>>>p0))&(&((~&(|$signed(p3))))));
  assign y9 = {1{{4{p8}}}};
  assign y10 = {(~(-{3{p11}})),{1{(|{3{p15}})}},(~&({2{p2}}=={1{p1}}))};
  assign y11 = (-{3{(4'd4)}});
  assign y12 = {2{{{2{b5}},{p0,p7,p9},(p15!=p16)}}};
  assign y13 = ({(a2<<<p3),(a2<<b3),{a2,p4}}<((a5&p8)&&(b3>=p2)));
  assign y14 = (((p5-p3)<<<(a5+b3))|((b3<b4)===(b0>b4)));
  assign y15 = (4'sd7);
  assign y16 = (((3'd3)>(b3!==b1))==($unsigned(((4'd8)<(b4!=a4)))));
  assign y17 = (~(a4^~a5));
endmodule
