module expression_00901(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-5'sd7);
  localparam [4:0] p1 = ((~|(5'd7))>>>((5'sd0)>>>(4'd2)));
  localparam [5:0] p2 = (3'd6);
  localparam signed [3:0] p3 = ({((3'd4)<=(3'd2)),((-4'sd7)<<(5'd14)),(+(-4'sd0))}===(((-3'sd1)!=(2'd3))^~((5'd4)!=(-4'sd4))));
  localparam signed [4:0] p4 = (~^(+((-2'sd1)!==((!((5'd3)>>>(5'd14)))^(~|(2'sd0))))));
  localparam signed [5:0] p5 = (-(^(&(((4'd7)===(3'd7))&(~&(4'd6))))));
  localparam [3:0] p6 = ((((4'd10)?(-3'sd3):(5'd26))>((2'sd0)?(3'd2):(4'd9)))^((3'd1)?(-3'sd1):(5'd8)));
  localparam [4:0] p7 = ((~&(~^(-{(2'sd0)})))>>((~(2'd3))&((2'd2)==(2'd2))));
  localparam [5:0] p8 = (((2'sd0)?(2'sd1):(5'sd7))?((4'd11)?(4'd14):(2'd0)):((5'd6)?(-4'sd2):(2'd3)));
  localparam signed [3:0] p9 = (((~^(4'd2))===((2'sd1)^(2'd3)))|({(2'sd0),(2'sd1),(2'd1)}>>((-4'sd6)?(2'd3):(4'd7))));
  localparam signed [4:0] p10 = {(-2'sd1),(-3'sd0),(5'd3)};
  localparam signed [5:0] p11 = (~^(4'd10));
  localparam [3:0] p12 = (({2{(5'd26)}}||{4{(2'd0)}})^(((-4'sd1)?(-3'sd2):(-4'sd6))?(4'd2 * (5'd27)):(3'd3)));
  localparam [4:0] p13 = (+(|{((3'sd0)|(5'd25))}));
  localparam [5:0] p14 = (4'd8);
  localparam signed [3:0] p15 = (|({(-4'sd3),(3'd3),(-2'sd0)}||(~(-5'sd12))));
  localparam signed [4:0] p16 = (^{3{((-2'sd0)?(4'sd7):(5'sd15))}});
  localparam signed [5:0] p17 = (!((-((2'sd1)>=(3'd4)))%(3'd0)));

  assign y0 = (~^(!(~&((&({p0,p1}&{{p5}}))||(-3'sd1)))));
  assign y1 = (~&(~|((p7?a2:a1)?(~^(|(b1?b3:p10))):((!b1)!=(b4|p15)))));
  assign y2 = (|(+(((!(-(b0^a4)))+(~^(a1?b2:b1)))===$signed(({{a1}}||({b4}))))));
  assign y3 = ((~^(~|(({3{p1}}<<<(&p3))>((a5!==a5)>(p10?p14:p7)))))+(^(~|(-({3{p10}}+(p14?p10:p12))))));
  assign y4 = (b0?a0:b5);
  assign y5 = {3{({2{a4}}?{3{b2}}:(a3?b1:b3))}};
  assign y6 = (!{((((a1^b0)-{a0,b4})==={a2,b4,a3})>>(((a3||b1)>(~|p14))>>(|(~(a5|a4)))))});
  assign y7 = (-(~|{4{{3{p15}}}}));
  assign y8 = (a3!==b2);
  assign y9 = (((&p1)<(a4||p1))==((~a5)&&(~&a4)));
  assign y10 = (~|((((a2==a5)^(+a2))!=(~&({4{a0}}!=(~&a3))))!==(~|{4{(~|b4)}})));
  assign y11 = {({b3,p6}?(b1<<b1):{4{p4}}),(((a2?a0:p13)?$signed(b5):{p6,p0})),(~^{(4'd2),{(a2&p8)}})};
  assign y12 = (((b0?a0:b5)===($signed(b0)-(-a5)))===({a0,b3,b2}?(^(b5<<<a4)):{a1,a0}));
  assign y13 = (~^(|($unsigned((^{((^(~a5))),{{3{a2}}},((-a3)>=(a0^a1))})))));
  assign y14 = ((4'sd4)&&((3'sd2)!=(a2%b1)));
  assign y15 = (~^{p14,p10});
  assign y16 = (&{({p0,b5,p9}<={a2,p11,p8})});
  assign y17 = (2'd3);
endmodule
