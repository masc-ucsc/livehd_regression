module expression_00433(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(!((5'd2 * (3'd7))/(-3'sd2))));
  localparam [4:0] p1 = {3{(~|{4{(3'sd2)}})}};
  localparam [5:0] p2 = (+(4'd13));
  localparam signed [3:0] p3 = {4{{2{(-2'sd1)}}}};
  localparam signed [4:0] p4 = (((((2'd0)<<<(-5'sd1))>=((3'sd2)==(2'd3)))<<<(((-4'sd4)||(3'd6))|((-3'sd2)*(2'd0))))<<((((4'd7)<=(4'd8))^~((-3'sd2)&&(5'd14)))>=(((3'sd3)/(4'd15))<<((2'd3)!==(2'sd0)))));
  localparam signed [5:0] p5 = ({((5'd4)<=(5'd12)),{(4'd6)},((5'sd9)!=(-2'sd1))}^~(((2'd2)^(-2'sd0))>((3'sd0)||(4'sd1))));
  localparam [3:0] p6 = (-5'sd9);
  localparam [4:0] p7 = (((-5'sd1)-(-3'sd2))-{(4'd13)});
  localparam [5:0] p8 = (~(-(-(((2'sd1)>>>(-3'sd0))==(&{(4'd12),(4'sd7)})))));
  localparam signed [3:0] p9 = ((5'd25)-(4'd3));
  localparam signed [4:0] p10 = (|(({(4'd6),(-5'sd12),(4'sd6)}<<<((-5'sd7)&&(3'd4)))^~(+((-5'sd3)==(3'sd1)))));
  localparam signed [5:0] p11 = {(({(-4'sd5),(-4'sd4)}<=((-2'sd1)&&(2'd2)))|((5'd2 * (5'd3))>>{(3'd1),(-2'sd1)}))};
  localparam [3:0] p12 = ((5'd13)?(2'd0):(4'd13));
  localparam [4:0] p13 = ((((5'sd14)^(5'sd12))?((-5'sd15)?(-5'sd0):(5'd4)):((-4'sd2)===(4'd15)))-(((4'd15)>>>(2'd2))%(-4'sd2)));
  localparam [5:0] p14 = {4{(4'd15)}};
  localparam signed [3:0] p15 = ((^({4{(2'd1)}}?{1{(4'd12)}}:((-4'sd4)?(5'd19):(5'sd11))))<{3{(|(3'd3))}});
  localparam signed [4:0] p16 = (~&(-(~|((^(-(-2'sd1)))?(~^(~^(5'd31))):((-5'sd13)?(2'd2):(-4'sd0))))));
  localparam signed [5:0] p17 = (({4{(-4'sd7)}}&&(5'd2 * (4'd7)))>>>({2{(-2'sd0)}}||{2{(4'd1)}}));

  assign y0 = (p4!=p16);
  assign y1 = (((b3?b2:a0)?(b1-b5):(a4!=a0))==={(b2?a2:b4),(b0>>b4),{a5,a1}});
  assign y2 = {1{{4{(a4?a5:b3)}}}};
  assign y3 = (p6&p0);
  assign y4 = (-((~&(p16>=p10))/p10));
  assign y5 = ((^{3{(2'd3)}})<<<({4{p17}}|(p9&b5)));
  assign y6 = (|($signed(a4)?(p4<<<a3):(~|p8)));
  assign y7 = {$signed(b5),{a3},{a2,a2}};
  assign y8 = $unsigned({{{p6,b1,a2},{p13,a4,a2}}});
  assign y9 = (2'sd1);
  assign y10 = (a4>p13);
  assign y11 = (((p8%p17)?(p1?p16:p4):(p10>=p7))||(((p7^~p2)>>>(p3?a2:p1))==(p6?p16:p1)));
  assign y12 = {2{$signed(({4{b2}}!=={3{a3}}))}};
  assign y13 = ({(((b1?b4:b5)<<<{p8})<$signed((b5?a4:a4)))}<((b2<p1)?{b2,b0,p2}:{2{p15}}));
  assign y14 = (({3{b2}}^~{(~^a5),{4{a4}}})!={(|(a2==a0)),{a4,p9,p4}});
  assign y15 = {{p12,b4},{p9,p0,p6}};
  assign y16 = (!(~&({2{b1}})));
  assign y17 = {3{(4'sd3)}};
endmodule
