module expression_00296(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{((4'sd7)!=(5'd10))},{{(-3'sd2),(2'sd1),(4'sd2)}}};
  localparam [4:0] p1 = ((~|{1{((-3'sd0)==(2'sd1))}})-(6'd2 * ((2'd0)>=(4'd9))));
  localparam [5:0] p2 = {(-{(|{(-(&{(-3'sd1),(4'd15),(3'sd1)}))})}),{{(2'sd1),(4'd11),(5'd28)},{(4'sd2),(3'd7)},(&{(-2'sd0)})}};
  localparam signed [3:0] p3 = (-4'sd4);
  localparam signed [4:0] p4 = (3'd0);
  localparam signed [5:0] p5 = (!({3{(3'd7)}}||(((5'sd12)===(3'd2))===((5'sd5)^(4'sd4)))));
  localparam [3:0] p6 = (((-3'sd0)<(-3'sd2))&&{3{(-4'sd6)}});
  localparam [4:0] p7 = ((4'd3)+(5'd2));
  localparam [5:0] p8 = {(3'sd1),(((3'sd3)===(5'sd10))>={(3'sd1),(5'd1)})};
  localparam signed [3:0] p9 = ((5'sd12)&((-3'sd2)===(4'sd6)));
  localparam signed [4:0] p10 = ((4'sd5)?(4'd15):(5'sd13));
  localparam signed [5:0] p11 = ({3{((4'd8)>(-5'sd11))}}!==({1{(-5'sd5)}}+{3{(3'd7)}}));
  localparam [3:0] p12 = ((-3'sd1)?(~(|((4'd2)>>>(2'd0)))):(~^(^(-3'sd2))));
  localparam [4:0] p13 = {{(-{2{{3{(-4'sd1)}}}}),((~|{(-4'sd2)})>>>(+(!(4'd7))))}};
  localparam [5:0] p14 = ((((-4'sd2)?(4'sd7):(3'd7))|((-4'sd3)>=(2'sd0)))!=(((3'd1)?(-3'sd2):(-5'sd4))-((-2'sd0)<(-4'sd7))));
  localparam signed [3:0] p15 = (2'd2);
  localparam signed [4:0] p16 = ({(5'sd2),(5'sd15),(2'sd0)}?(~^((3'sd3)>>>(-4'sd0))):(|(!(4'd8))));
  localparam signed [5:0] p17 = ({1{{3{(2'sd0)}}}}?({1{(3'd4)}}?((2'sd0)&&(2'sd1)):(^(-5'sd11))):(((3'd1)?(5'd10):(3'sd0))?((-3'sd2)||(4'd15)):((4'd11)>(2'd3))));

  assign y0 = (5'sd7);
  assign y1 = ((2'sd1)?(5'd2 * (5'd24)):((2'sd1)));
  assign y2 = (5'd27);
  assign y3 = (~^(((p5?p11:a0)?(p9?a3:b1):(^(p6?p6:p4)))|((a5===a5)%b3)));
  assign y4 = ((b5==b5)!==(b5!=a5));
  assign y5 = (~|(~(~|(5'd11))));
  assign y6 = (|a4);
  assign y7 = {3{(|(a2<<b0))}};
  assign y8 = ((p0?p7:p12)?(p4^~b2):(b2?p16:b2));
  assign y9 = (~^(~&(({2{b4}}!==(~&b1))!==(!{4{b3}}))));
  assign y10 = $signed((a5?b0:b5));
  assign y11 = ((4'd2 * (!(6'd2 * p2)))+((p16<p12)^(b5!==b2)));
  assign y12 = (~|(-(({a3,b0}||(-{a4}))-(-({b0,a5,b4}-(~|b5))))));
  assign y13 = (~(-3'sd3));
  assign y14 = (((b5+b2)<<(+b2))!==({b0,a0,a1}<<<{b2,b0}));
  assign y15 = (((a3?a1:b5)?$unsigned(b1):(+a2))||((a4%a0)>=(~(p16<=a4))));
  assign y16 = (~^(&{2{b3}}));
  assign y17 = (~|(&(+(4'd2))));
endmodule
