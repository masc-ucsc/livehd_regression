module expression_00803(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{{2{(5'd24)}}}};
  localparam [4:0] p1 = {(|(4'd2 * ((4'd15)==(5'd22)))),(((3'd1)==(4'sd2))?((3'd7)?(2'd1):(3'sd0)):((5'd14)?(-3'sd2):(-3'sd1))),(-(((-3'sd2)!=(-4'sd1))|((5'd17)>=(5'sd11))))};
  localparam [5:0] p2 = {3{(3'sd1)}};
  localparam signed [3:0] p3 = ((-5'sd10)^(2'd3));
  localparam signed [4:0] p4 = {({((3'd0)^(3'd6))}?((2'd3)==((2'd3)?(2'd1):(-5'sd15))):((3'd3)?(5'd22):(5'd0)))};
  localparam signed [5:0] p5 = {(((3'sd3)>>>(-4'sd3))?(-5'sd11):{(-2'sd0)}),(3'sd2)};
  localparam [3:0] p6 = ((3'sd1)?(4'd0):(4'd6));
  localparam [4:0] p7 = {1{(4'd7)}};
  localparam [5:0] p8 = {(^(~|(~^(-4'sd0))))};
  localparam signed [3:0] p9 = ((((4'd6)?(-5'sd1):(-2'sd0))===(-(2'd1)))>(^(|((5'd12)>(5'd30)))));
  localparam signed [4:0] p10 = ((((2'd2)^~(-5'sd6))>=(!(4'd5)))<<<((~(4'sd7))||((-4'sd4)<(3'd6))));
  localparam signed [5:0] p11 = (!{2{(!(&(&((5'sd13)?(3'd6):(3'd4)))))}});
  localparam [3:0] p12 = ((4'd11)^(5'd25));
  localparam [4:0] p13 = {{4{(-4'sd2)}}};
  localparam [5:0] p14 = {3{((5'd29)?(2'd2):(5'sd5))}};
  localparam signed [3:0] p15 = {2{(5'd3)}};
  localparam signed [4:0] p16 = ({1{((2'sd1)+(-3'sd2))}}?((3'sd0)>(2'd3)):{1{((-2'sd1)|(4'd5))}});
  localparam signed [5:0] p17 = ((((-5'sd14)<(2'd1))<<((-3'sd2)>=(4'd14)))-(((5'd13)^(2'd0))>>>{(3'd3),(2'd3)}));

  assign y0 = ((p16|p2)^{4{p13}});
  assign y1 = {1{{2{(~(~{1{p2}}))}}}};
  assign y2 = {(~&(-(!((b1&p14)<<<(a4^~p16))))),(~^{(~|((b5!=p6)&&(p14&&p2)))})};
  assign y3 = (!(&{({(p2?p12:b1),(p9?p16:b2)}?{{a5,a0},{4{a3}}}:{2{(b4^a3)}})}));
  assign y4 = {4{{{2{p9}}}}};
  assign y5 = (b5+b5);
  assign y6 = ({3{(a5===a2)}}+({4{a0}}<{p7,b1}));
  assign y7 = ((((p14?p17:p14)?(b1?b1:p2):(p7?b2:p5))&((p12>>>p7)>>>(p2^p3)))<=({1{{b1,p13}}}?(a2==p11):{(b2?p2:p8)}));
  assign y8 = $unsigned((({1{{(((3'sd3)<<<{(-4'sd3)})>{3{(a1-b3)}})}}})));
  assign y9 = {{a2,a3},((3'sd1)),(|(p4<a1))};
  assign y10 = (((b0&b0)*(p11+b1))!=((a2^~b0)%p17));
  assign y11 = (^$unsigned(({{2{b4}},{2{a4}}}+(!{(~|p14)}))));
  assign y12 = (&(((a5&a3)<<<(a5>=b3))==((6'd2 * b0)?(~&p6):(p16-a4))));
  assign y13 = (~^(((|(a2!==a2))!=(~(a3<<<b4)))^~(-((a5|a2)===(|(|b3))))));
  assign y14 = (5'd2 * $unsigned((p8?a1:a4)));
  assign y15 = (({p11,a3,p7}?(5'd11):(-3'sd1)));
  assign y16 = ((p11<<<p11)?(a3?a2:p12):(a1%p5));
  assign y17 = (((~^(~&p17))<(&(~&p16)))|(~((^(~^(^(p9==p14)))))));
endmodule
