module expression_00077(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd9)?(-3'sd3):(2'd0))>(+((5'd5)?(4'sd6):(2'd2))));
  localparam [4:0] p1 = ({(((-5'sd9)&(-5'sd14))?{(-5'sd14)}:((2'd3)?(5'd7):(3'sd3)))}!=(4'd12));
  localparam [5:0] p2 = (~&(^{2{(~|{1{(&(~&(~(-4'sd6))))}})}}));
  localparam signed [3:0] p3 = ((4'd3)||(2'd2));
  localparam signed [4:0] p4 = ({(4'sd5),(-4'sd7)}?((5'd8)^~(3'd6)):((2'd3)<<(3'd6)));
  localparam signed [5:0] p5 = (!{1{{4{(|(2'd0))}}}});
  localparam [3:0] p6 = (-4'sd4);
  localparam [4:0] p7 = (((5'd3)?(3'sd0):(4'd7))^~((4'd2)?(2'd2):(2'd3)));
  localparam [5:0] p8 = (5'd16);
  localparam signed [3:0] p9 = ((5'd2)+(((5'sd7)<(4'sd2))&&(3'd6)));
  localparam signed [4:0] p10 = (~&(-4'sd1));
  localparam signed [5:0] p11 = (-{4{(5'sd3)}});
  localparam [3:0] p12 = (4'd5);
  localparam [4:0] p13 = (&((4'd15)^(~^{2{(|((5'sd5)!==(3'd7)))}})));
  localparam [5:0] p14 = ((~^(5'd6))?(!(6'd2 * {2{(4'd6)}})):(((5'd1)==(4'd15))-(~^(3'd2))));
  localparam signed [3:0] p15 = ((!((3'd0)?(2'sd1):(5'd15)))?(~|((5'd2)?(2'd2):(3'd7))):((~|(5'sd13))?((5'sd4)?(-2'sd0):(4'd12)):(^(-5'sd6))));
  localparam signed [4:0] p16 = (-3'sd2);
  localparam signed [5:0] p17 = (((-2'sd1)^~(5'd3))%(5'd4));

  assign y0 = {3{(|(b1-b5))}};
  assign y1 = (~&$unsigned((b2!==a3)));
  assign y2 = ($signed(p4)?(p3):(p0==p1));
  assign y3 = (((3'sd2)!==(-5'sd9))|(((5'sd4)<(3'sd3))<<(2'd0)));
  assign y4 = ($signed(({1{a5}}&{2{b3}})));
  assign y5 = ((a5==b1)?(-3'sd1):(p6|p1));
  assign y6 = $signed({{$signed(a5),(~p14)},{$signed({b5})},(^(a1===b4))});
  assign y7 = (&(({(p5||p9),(~&(&p16))}?((p13?p3:b3)!={$signed(p10)}):(-{4{b2}}))));
  assign y8 = (-2'sd0);
  assign y9 = $unsigned((~|(5'd3)));
  assign y10 = ((((b5&b1)==(b1^b4))<=((a2|b2)^~(b1<b1)))!==(((|b1)!==(+a2))>((~^b5)<(b4-a4))));
  assign y11 = ((-(!(5'sd11)))&&(~|(-5'sd0)));
  assign y12 = (((a5!=p8)!=(a5?b5:a1))|((2'sd0)+(a5!=p7)));
  assign y13 = {(-(p1?p4:p13))};
  assign y14 = {3{(^(^{1{{3{a3}}}}))}};
  assign y15 = (!(|p3));
  assign y16 = (~&{3{a3}});
  assign y17 = {(^{{3{a1}},{2{a0}},{1{b2}}}),(+(~(&(-(a3>>b4)))))};
endmodule
