module expression_00964(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-4'sd0)>>(5'sd14))||(~&(-2'sd1)));
  localparam [4:0] p1 = (|(^(-({{(5'sd4),(2'd3)},((4'sd6)^~(4'd14)),{(3'd3),(-5'sd5),(5'sd1)}}>>(^(+{(5'sd9),(-2'sd1),(4'd3)}))))));
  localparam [5:0] p2 = (|(((2'd1)!==(-4'sd2))|(+(2'd1))));
  localparam signed [3:0] p3 = (-5'sd11);
  localparam signed [4:0] p4 = ((-((3'd4)&(3'd7)))%(4'sd6));
  localparam signed [5:0] p5 = ((4'sd2)!==(4'd5));
  localparam [3:0] p6 = (!({1{(3'd2)}}?(((-3'sd3)?(5'd21):(3'd1))&{1{(2'sd1)}}):{2{{2{(3'sd2)}}}}));
  localparam [4:0] p7 = (((5'd8)^~(4'd13))!==((2'sd0)<(-4'sd3)));
  localparam [5:0] p8 = (&(((5'd9)>>>(2'd2))===((5'd20)|(4'd15))));
  localparam signed [3:0] p9 = (((-5'sd14)?(~(3'sd2)):(6'd2 * (2'd0)))?(^(~|(4'd8))):{((4'd9)&(5'd2)),(!(-5'sd11)),(!(2'sd1))});
  localparam signed [4:0] p10 = (!(-((-2'sd1)>>(-4'sd1))));
  localparam signed [5:0] p11 = (~^(4'sd6));
  localparam [3:0] p12 = {4{(2'd2)}};
  localparam [4:0] p13 = {(+(-{(3'd0),(-4'sd3),(-4'sd4)})),{(5'd22),(2'sd1),(-3'sd0)},{{(3'd2)},{(5'd1),(4'sd7),(4'sd0)}}};
  localparam [5:0] p14 = (~((~|{(^(2'sd0)),((-5'sd0)<<<(5'd14))})^{{((4'd8)?(-5'sd11):(2'd0))}}));
  localparam signed [3:0] p15 = ({2{(-5'sd14)}}?{1{(-2'sd0)}}:((5'sd4)?(2'd2):(-3'sd1)));
  localparam signed [4:0] p16 = ((((2'd3)!=(4'd9))?((5'sd13)<<(2'sd1)):((5'sd6)?(5'd12):(4'd14)))+((2'd1)<<((5'd22)?(-2'sd1):(2'd0))));
  localparam signed [5:0] p17 = {(4'd2 * (&(4'd15))),((4'sd3)?(4'sd7):(4'd6)),{(~&(3'd0)),((-5'sd14)>>>(4'sd2))}};

  assign y0 = (~&(((5'd2 * (p2||b2))^~((a0>a1)|$unsigned(a1)))-(((a2!=b3))===(5'sd1))));
  assign y1 = (p0<<<p8);
  assign y2 = {{{1{{3{{4{p7}}}}}}}};
  assign y3 = (((a3?a4:b2)?(a2?b4:a2):(b1?b0:a3))?((b5?a3:p10)?(b3?b3:b0):(a5?a0:b5)):((b5?b1:b4)?(a4?p10:b4):(a5?b4:b5)));
  assign y4 = (3'd3);
  assign y5 = ((p15==p12)/p2);
  assign y6 = (((b3>>>a3)?(a4===a1):(a4))?((a3?a1:b1)&&{b3,b4}):($signed(b1)?(-b5):(-a4)));
  assign y7 = (({3{a5}}?(a5):{a3})?{4{b4}}:(4'd5));
  assign y8 = (~&(|((-((&(a0===a3))>=(+(~b0))))-(^(3'd5)))));
  assign y9 = (!(-3'sd2));
  assign y10 = (~^(-2'sd0));
  assign y11 = ((+(~(-(~&p6)))));
  assign y12 = (6'd2 * {p6,p2,p14});
  assign y13 = ((((5'd5)>>>(4'd1))+((a4>a3)%a3))==(-5'sd12));
  assign y14 = (2'd1);
  assign y15 = {a2,a1,p9};
  assign y16 = (2'd1);
  assign y17 = (-$unsigned({{({{$signed((-b4))},(b1?a2:a0),(b1?a0:p4)})}}));
endmodule
