module expression_00172(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^{(4'sd1),(4'sd6),(5'd6)});
  localparam [4:0] p1 = {(6'd2 * (2'd0)),{(2'd3)}};
  localparam [5:0] p2 = (!(2'd2));
  localparam signed [3:0] p3 = (|(~((~&(3'd3))>>>((4'sd7)||(2'd2)))));
  localparam signed [4:0] p4 = {(((-2'sd1)!=(-2'sd0))==={3{(4'd6)}}),{4{{2{(-2'sd1)}}}}};
  localparam signed [5:0] p5 = (+(+({{(-(5'd2)),{(5'd11)}}}!=(+(4'd2 * (5'd20))))));
  localparam [3:0] p6 = (5'd2 * (3'd0));
  localparam [4:0] p7 = ((5'd21)>>(5'd8));
  localparam [5:0] p8 = ((4'sd4)>(4'd2));
  localparam signed [3:0] p9 = (|((-(~|(&(~^((3'sd1)==(5'd2))))))>>((|((5'd10)<=(2'd1)))|(&(^(5'sd15))))));
  localparam signed [4:0] p10 = {2{(4'sd6)}};
  localparam signed [5:0] p11 = (~&(3'sd2));
  localparam [3:0] p12 = (3'd0);
  localparam [4:0] p13 = ((((2'd0)?(3'd3):(3'sd2))-(~|(5'sd5)))?{1{(((3'd2)?(3'sd3):(4'd13))!=={(5'd23),(5'sd4)})}}:(&{4{(4'd11)}}));
  localparam [5:0] p14 = {{((3'sd2)==(3'sd1))},(((-5'sd3)^~(2'd1))>=((3'd3)!==(-4'sd3))),(((4'd11)>>(-5'sd4))==((-5'sd11)^~(-4'sd3)))};
  localparam signed [3:0] p15 = {(&{1{{{4{(3'd5)}}}}}),(!(~&{2{(^{(4'd6),(5'sd6),(-3'sd1)})}}))};
  localparam signed [4:0] p16 = ((4'd2 * (4'd13))>=(-5'sd9));
  localparam signed [5:0] p17 = (5'd2 * ((4'd3)<=(2'd3)));

  assign y0 = (($unsigned(b0)||{2{b4}})?(-4'sd6):((p10)&(b0==b1)));
  assign y1 = (a1?a4:a2);
  assign y2 = (&{3{(~^(-{3{b2}}))}});
  assign y3 = (3'd5);
  assign y4 = {($signed((2'sd0))>((p17)?(b2?a1:p17):(p12>=b4)))};
  assign y5 = ((p0%p13)/p11);
  assign y6 = ((p8&p2)-(~&{2{p7}}));
  assign y7 = ((~&(4'd8))<<<(+(^(2'sd1))));
  assign y8 = ((4'd11)!=(p5||p2));
  assign y9 = {({{a0},(p3?b4:b1),(!b3)}<<<$signed((^((a4^~b5)!==(!b4)))))};
  assign y10 = (-{(((p12)==(a0<<<p2))&&{3{a5}}),(((a0||b0)!=={b1,b3,b0})=={b4,b0,a3})});
  assign y11 = ({1{(p8&b0)}}&{1{$unsigned((p10-p17))}});
  assign y12 = ({({b4,b5,a3}===(4'd14))}+(4'd2 * {p13,b2,p0}));
  assign y13 = $signed(({3{{4{b0}}}}^~{(~&b5),(a3)}));
  assign y14 = {1{{2{{4{b5}}}}}};
  assign y15 = {3{(a5)}};
  assign y16 = ((p15?p5:p13)?(4'sd2):(b2==b5));
  assign y17 = {(5'd8),$signed($signed(p13)),(~^{p10,a5,p15})};
endmodule
