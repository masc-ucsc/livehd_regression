module expression_00498(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(2'd3));
  localparam [4:0] p1 = ((((-5'sd2)|(-2'sd0))|{(5'd24),(3'sd0)})==(3'd1));
  localparam [5:0] p2 = (~&(5'sd5));
  localparam signed [3:0] p3 = (4'sd7);
  localparam signed [4:0] p4 = ((((4'sd4)/(2'sd1))<=((4'd5)>=(-2'sd0)))>=(((5'sd12)|(-2'sd0))^~((-2'sd0)||(2'd3))));
  localparam signed [5:0] p5 = (~^{4{(3'd1)}});
  localparam [3:0] p6 = ((((5'd28)!==(-3'sd1))^(&(2'd3)))>=(&(-(!((5'sd14)&(3'sd3))))));
  localparam [4:0] p7 = ((3'd4)?(2'd0):((3'sd2)?(-4'sd3):(4'd10)));
  localparam [5:0] p8 = (((-5'sd8)||(4'sd0))&{(4'd0),(5'd26),(4'd14)});
  localparam signed [3:0] p9 = (((2'd2)!==(3'd6))-(~&((2'd3)<<<(4'd11))));
  localparam signed [4:0] p10 = ((5'd11)?(2'sd0):(2'd0));
  localparam signed [5:0] p11 = (~|(&{{(-3'sd3),(2'd1),(3'd2)},((^(-3'sd2))>>{(3'd2)}),(!(5'd31))}));
  localparam [3:0] p12 = (4'd2 * ((4'd11)<(2'd1)));
  localparam [4:0] p13 = {{4{{(-2'sd1),(4'd11)}}},(!({4{(-4'sd5)}}<<(&(!(-3'sd3)))))};
  localparam [5:0] p14 = {(|((3'd2)<=(-2'sd1))),((4'd1)-(2'd0))};
  localparam signed [3:0] p15 = (~&((-4'sd0)<=(((-3'sd2)^(4'd8))===((-3'sd0)&(3'd5)))));
  localparam signed [4:0] p16 = (~&({{3{(4'sd0)}},((-3'sd1)<(2'd2))}?(|(~&(^((3'd2)==(5'd7))))):(((-5'sd7)?(-3'sd2):(-5'sd4))?{3{(5'd25)}}:{(3'sd2)})));
  localparam signed [5:0] p17 = ((((2'd1)>(5'sd8))>=((2'd1)===(-3'sd3)))==(~|(((4'd11)<<(3'd5))<=((3'sd1)>(4'd6)))));

  assign y0 = (5'd2 * b2);
  assign y1 = {(b2?p11:p3),(p11<p7),(p7^a0)};
  assign y2 = (&{{(6'd2 * (b1-p14)),((b3?a0:b4)&{3{b1}}),(6'd2 * (4'd11))}});
  assign y3 = {2{((b0!==b4)?(a4>a4):(b1|b0))}};
  assign y4 = (~&($unsigned({{$signed(p5)},(!(4'd10))})));
  assign y5 = ((+(^((!(2'd0))!=(p0&p12))))&&(4'sd2));
  assign y6 = (+(~|$unsigned((^(({1{{4{(a1>>a0)}}}}!==(((a3>>a5))===(^$unsigned(b4)))))))));
  assign y7 = ((b2<a4)?(!p11):{a3});
  assign y8 = (2'd0);
  assign y9 = {(((a4?b2:p8)>{(b3-b4),{p11}})<<<{(p6?a3:a1),(a0!==b1),(a3!==a2)})};
  assign y10 = (p4|a1);
  assign y11 = {4{(p10||a3)}};
  assign y12 = {(~|(((b4>>p4)&(4'd4))?{(a3?p3:p1),{a0},(2'd3)}:((2'sd1)||(3'd2))))};
  assign y13 = ((p1?p5:b5)?({2{a2}}>=(b1?b1:b4)):{p14,p5,a3});
  assign y14 = (-((a3-p16)<=(-4'sd0)));
  assign y15 = {p0,p10,a4};
  assign y16 = (p3?p15:a0);
  assign y17 = (&p7);
endmodule
