module expression_00040(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd8);
  localparam [4:0] p1 = ((3'd5)%(2'd0));
  localparam [5:0] p2 = {(2'd3),(-5'sd11)};
  localparam signed [3:0] p3 = (^{(&{(-5'sd5),((3'd3)<=(2'sd0)),((4'd5)<=(5'd8))}),(&{{(5'd4),(4'd13)},(2'sd1)})});
  localparam signed [4:0] p4 = (3'd7);
  localparam signed [5:0] p5 = (|((+(+{(-4'sd2)}))&{(5'd2),(5'sd8),(4'd1)}));
  localparam [3:0] p6 = (2'd2);
  localparam [4:0] p7 = ((((4'sd5)>>>(2'd2))!=(4'sd1))|(((-2'sd1)^~(-4'sd0))>((-4'sd0)%(-2'sd0))));
  localparam [5:0] p8 = ((((3'd4)==(2'sd1))^(^(3'd6)))>>(((-2'sd1)===(5'sd0))&&{4{(5'sd4)}}));
  localparam signed [3:0] p9 = (^(-5'sd1));
  localparam signed [4:0] p10 = ({2{{3{(5'sd3)}}}}>>(|(((-2'sd1)&&(3'd0))!==(5'd2 * (2'd3)))));
  localparam signed [5:0] p11 = (|((((4'sd0)<=(2'd1))^{(2'sd1),(2'd3),(4'd0)})?((~&(3'sd1))^((-5'sd14)&(-5'sd7))):(~(4'd2 * (5'd27)))));
  localparam [3:0] p12 = ((((-2'sd0)>=(-4'sd4))<=((-5'sd6)^(4'd13)))===(((3'd0)!=(3'd6))>>(5'd2 * (2'd0))));
  localparam [4:0] p13 = ((5'd8)>(5'sd15));
  localparam [5:0] p14 = ((~|(4'd3))?((3'd5)<<(-5'sd1)):((4'sd3)&&(5'sd10)));
  localparam signed [3:0] p15 = ((-((4'sd0)&&(5'sd13)))<<((5'd30)?(5'sd4):(2'sd0)));
  localparam signed [4:0] p16 = ({3{(5'd28)}}?(~|((4'sd0)>>(-2'sd1))):(((3'sd1)<<(2'd0))<=((4'd13)||(2'sd0))));
  localparam signed [5:0] p17 = {(-4'sd1)};

  assign y0 = (2'd1);
  assign y1 = (a1>>b3);
  assign y2 = ({4{(&p13)}}>{1{(+({1{a2}}?(p7?p12:p8):(-p4)))}});
  assign y3 = ((3'd2)>>>(4'd0));
  assign y4 = {1{{4{(4'd7)}}}};
  assign y5 = {{1{{4{(+b2)}}}},{(-(+(-3'sd1))),(4'sd4)}};
  assign y6 = {{{(~^(+{{{a1,b2,a4}},(&(b3&&a0)),(~^(!a1))}))}}};
  assign y7 = (~(~{2{p3}}));
  assign y8 = (p17>=b2);
  assign y9 = (-(((&$signed($unsigned($signed((!p5))))))>=$signed(((-(p7&p6))<(p7<b4)))));
  assign y10 = ({1{((^(p10<<p5))<((~&p11)-(~^p9)))}}||{2{({3{p5}}&(p2>=p9))}});
  assign y11 = (~^(~|(~&(~{(5'sd15)}))));
  assign y12 = ((~((|$signed(($signed($signed(a0))^(b1?p12:p6))))^(($signed((&$signed($signed($signed((p12?b4:p1)))))))))));
  assign y13 = (+(|((-4'sd3))));
  assign y14 = {({{{a0,a3},(+{a5,a4})}}===(^((-{b5,a2,b5})>>(a0<a2))))};
  assign y15 = ({p8}?(4'd2 * p2):(b4?p7:p8));
  assign y16 = ({b5,p0,p7}+(b0?p10:a5));
  assign y17 = (!$signed((((p11)^(a1<<p9))>>{2{(~^a2)}})));
endmodule
