module expression_00119(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(2'sd1)}};
  localparam [4:0] p1 = {2{(5'sd11)}};
  localparam [5:0] p2 = (({(3'd2),(5'd30)}>{{(3'd3)}})+{(((2'd0)-(4'd8))>>((-2'sd1)<<<(4'sd5)))});
  localparam signed [3:0] p3 = ((-5'sd13)?(5'd13):(4'd10));
  localparam signed [4:0] p4 = ((4'd3)?(5'd24):(-2'sd0));
  localparam signed [5:0] p5 = {1{({2{(2'sd0)}}?{(5'd31)}:{1{(-5'sd4)}})}};
  localparam [3:0] p6 = {1{(3'sd0)}};
  localparam [4:0] p7 = ((4'd8)>>(4'sd5));
  localparam [5:0] p8 = (&(~((-4'sd7)<<<(+(((3'd1)>=(3'd6))?((-3'sd0)-(5'sd15)):(-(5'd27)))))));
  localparam signed [3:0] p9 = ((5'sd1)>>>(-5'sd3));
  localparam signed [4:0] p10 = (((2'd3)&((2'd3)==(-3'sd0)))^(((5'd16)|(2'sd0))!=((5'd18)/(5'd6))));
  localparam signed [5:0] p11 = (((2'd0)?(4'd14):(2'd3))^((2'd0)||(3'd6)));
  localparam [3:0] p12 = (~|(~((((3'sd3)^~(3'sd3))<=(~|(-(2'sd0))))<<<(((3'sd3)<<<(2'sd0))?(|(-2'sd1)):((5'd13)?(5'd14):(5'd16))))));
  localparam [4:0] p13 = (5'd2 * (~&(~^(2'd1))));
  localparam [5:0] p14 = (~^((((-5'sd9)?(3'd5):(3'd2))<=(~(-4'sd3)))?{((-5'sd15)^~(2'd0)),((4'd6)<<(-4'sd6))}:((~^(2'sd1))+(|(-2'sd0)))));
  localparam signed [3:0] p15 = (&((2'd1)?(3'd7):(5'sd6)));
  localparam signed [4:0] p16 = ((-5'sd7)%(3'sd1));
  localparam signed [5:0] p17 = (((5'sd12)&(+(4'd3)))>=(2'd0));

  assign y0 = (p4<p13);
  assign y1 = ({(|p14),(p2<<<a5)}>(~|(&{p12,p2})));
  assign y2 = (~((p14)<<<{p10,a2}));
  assign y3 = (~(!$signed(p1)));
  assign y4 = ((3'd3));
  assign y5 = $unsigned((((4'sd5)<$signed($signed((($signed((-3'sd0))||(3'd7))))))));
  assign y6 = (!((p11!=p5)<<(p6>p16)));
  assign y7 = $unsigned(b3);
  assign y8 = (3'd1);
  assign y9 = (-3'sd1);
  assign y10 = (((b3?p14:a3)+(p0?a5:a5))?($unsigned(p11)?$unsigned(b2):$unsigned(a4)):$signed(($unsigned(b1)|{1{b4}})));
  assign y11 = (4'sd0);
  assign y12 = (-4'sd2);
  assign y13 = (-5'sd2);
  assign y14 = $unsigned({4{p8}});
  assign y15 = ({(a0!=a2),(b0===b0)}===(~^({a1,a3,a1}<(b4>=b4))));
  assign y16 = {{({2{p11}}-{3{p0}})},(3'sd1)};
  assign y17 = (~(-2'sd1));
endmodule
