module expression_00988(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{((-2'sd1)>((-5'sd7)>>>(3'd4)))}};
  localparam [4:0] p1 = {4{(3'sd1)}};
  localparam [5:0] p2 = (((~(3'd3))>>((-3'sd3)?(-2'sd1):(4'sd4)))||((|(5'd11))%(2'd3)));
  localparam signed [3:0] p3 = (-5'sd7);
  localparam signed [4:0] p4 = (((-4'sd6)&(-5'sd3))+((3'd7)!=(4'sd0)));
  localparam signed [5:0] p5 = (~|(^{{(4'd9),(2'd1),(4'd10)},{1{{(2'sd1)}}}}));
  localparam [3:0] p6 = {{2{(~(3'sd1))}}};
  localparam [4:0] p7 = ((-(-3'sd2))===(3'sd2));
  localparam [5:0] p8 = (~^((~(~|(((5'sd10)^~(-5'sd15))?(~&(4'd11)):{2{(-4'sd7)}})))^(((3'd3)?(2'sd1):(3'sd2))<<{2{(4'd10)}})));
  localparam signed [3:0] p9 = {((~^(~&((4'sd7)+(3'sd0))))<=((4'sd3)<<((3'sd2)===(4'sd1))))};
  localparam signed [4:0] p10 = {2{(5'd12)}};
  localparam signed [5:0] p11 = ((5'd15)|(5'sd13));
  localparam [3:0] p12 = ((-3'sd0)?(3'sd3):(-4'sd1));
  localparam [4:0] p13 = ((((5'd10)!=(-3'sd1))-((3'sd2)<<<(4'sd7)))&&(5'd2 * ((2'd1)!==(5'd1))));
  localparam [5:0] p14 = ((+((5'sd10)>>(2'sd0)))>>((2'd2)^(4'd8)));
  localparam signed [3:0] p15 = (|{3{(+(-4'sd4))}});
  localparam signed [4:0] p16 = (5'sd8);
  localparam signed [5:0] p17 = {1{(~^{4{((4'sd3)^(2'sd1))}})}};

  assign y0 = {(~|(+(~|(!(6'd2 * (+b2)))))),((^(p10-b3))?(!(p5||b4)):(b2>>>p8))};
  assign y1 = (&(a4<<<p9));
  assign y2 = (&(+(!(&(~&((~|(|(~p14)))))))));
  assign y3 = (-{(|{(~&(!b5)),(~&{p12,p6})}),{4{(p3)}}});
  assign y4 = (((2'd3)&(-4'sd4))!==((5'd2 * (a1<<a2))!==(2'sd0)));
  assign y5 = {4{{p12,p2,p8}}};
  assign y6 = (~&{{{b4,a5}}});
  assign y7 = ((^((b4>p6)?(p2>>p16):(-4'sd4)))&&(|((p9>>a5)*(p8?p3:b5))));
  assign y8 = (~|((3'd7)?(-3'sd3):{{4{b3}}}));
  assign y9 = {3{{{2{p12}},(3'd6),(5'd2 * p7)}}};
  assign y10 = (({1{($unsigned(p16))}}>>>(+(+(p16))))>>(+{3{(p10>>b0)}}));
  assign y11 = (^{4{{p8,p17}}});
  assign y12 = (5'd6);
  assign y13 = (~^(~&(~|(~|(~^(~^(4'd2 * (-(~&b0)))))))));
  assign y14 = {(~^{(3'sd2)})};
  assign y15 = {1{((b3?b1:a0)&&((+a1)==(~|b5)))}};
  assign y16 = {4{{2{(p3?p2:p13)}}}};
  assign y17 = ((|{2{(b4<b0)}})&($signed((b4^~p13))>$unsigned((+p16))));
endmodule
