module expression_00900(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((5'd18)^(2'd1))>=((4'sd1)*(4'd1)))?((5'd8)===((3'sd0)&&(3'd7))):(((3'd5)?(-5'sd2):(3'd3))||((4'd9)?(3'd4):(2'd0))));
  localparam [4:0] p1 = (((4'd3)<(-5'sd10))<=((4'd10)^(-2'sd1)));
  localparam [5:0] p2 = (((3'sd2)<=(5'd10))-(|{(5'd25)}));
  localparam signed [3:0] p3 = (((2'd1)>>(5'd18))/(2'd1));
  localparam signed [4:0] p4 = (|(((4'd2)?(-3'sd2):(3'd2))?((3'd4)?(5'sd2):(3'd4)):(-((-2'sd1)?(5'd16):(2'sd1)))));
  localparam signed [5:0] p5 = ((((4'sd6)>=(2'd2))+((2'sd1)<(2'd3)))&&(((3'sd0)==(-3'sd1))&((5'd0)<(4'd10))));
  localparam [3:0] p6 = ({3{(4'd6)}}+{2{{(3'd0),(3'd2),(-5'sd5)}}});
  localparam [4:0] p7 = {(-2'sd0),(-2'sd1)};
  localparam [5:0] p8 = (5'd26);
  localparam signed [3:0] p9 = ((-2'sd1)<<<(-2'sd1));
  localparam signed [4:0] p10 = (~&((~^(((4'd2)/(-3'sd2))&&((4'sd4)?(2'd3):(2'd2))))?(((-4'sd1)==(4'sd2))>>>((5'd15)?(-2'sd1):(-5'sd8))):((!(4'd3))+((-4'sd4)-(5'sd2)))));
  localparam signed [5:0] p11 = ((-4'sd7)?(-2'sd1):(-4'sd6));
  localparam [3:0] p12 = (((5'd16)==(2'sd0))?((-5'sd0)?(2'd0):(2'd3)):((4'd11)>=(4'd4)));
  localparam [4:0] p13 = (!(-(~^(6'd2 * (^(~&(2'd0)))))));
  localparam [5:0] p14 = ((3'd2)+(4'sd2));
  localparam signed [3:0] p15 = (!(&{4{(2'd2)}}));
  localparam signed [4:0] p16 = (~^((~^(+(~|{(4'd6),(2'd0),(4'd1)})))==((~|(4'sd0))>>{(3'd1),(3'sd2),(-2'sd1)})));
  localparam signed [5:0] p17 = ((+(-2'sd0))<<<((-4'sd4)&(4'd5)));

  assign y0 = ({((-a3)?(b5?b5:p8):{4{a2}})}?({b4}?{a4,b2,b2}:(b5?b3:b1)):(^{(&b2),(-a2),{2{a3}}}));
  assign y1 = (2'd2);
  assign y2 = (!(~^((+((a1===b3)?(|p16):(p8>>p15)))<<<((+(b0!==b2))?(p8?p14:p14):(p9>>>b3)))));
  assign y3 = {2{(|{2{b4}})}};
  assign y4 = (4'sd4);
  assign y5 = (|(((4'd2 * (a2^~a2))<={1{(b4>>>b4)}})^((!(+(b5&a2)))<=((a0==a2)>=(b0!==a2)))));
  assign y6 = {(|(~&{4{{p9,p4,p6}}})),(^{4{{1{p13}}}})};
  assign y7 = (((5'sd6)<(-2'sd0))==(~(~^(!{4{b4}}))));
  assign y8 = (^({{p12,a0,p3},(&p12),(p11<p9)}>>(~&(2'd0))));
  assign y9 = {4{{3{p17}}}};
  assign y10 = (((a2&&b1)<=(b2==a3))?((b2>>p16)&(b2?b2:b2)):{((p4))});
  assign y11 = ($signed((b4-b4))<=(p0==p4));
  assign y12 = (~((~^(^(4'd3)))^((b1>=a1)==(5'd23))));
  assign y13 = ((~&(&(~|{p16,p17})))<(|(|(~&(p17+p17)))));
  assign y14 = (5'd26);
  assign y15 = (-3'sd1);
  assign y16 = (((b5|b5)^~(-{a1,a3,b3}))?((b1?b1:a0)<<<{(b3+b1)}):({b1}?{a4,b1}:(b3|a1)));
  assign y17 = (~((~|((((~&p11)<=$unsigned(a5)))))&(~&((~$signed(b3))-(+(b0<a2))))));
endmodule
