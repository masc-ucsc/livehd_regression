module expression_00357(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd13)&&(5'd5))&((3'd3)===(4'sd0)))>>>(((5'd11)!==(5'd2))!==((5'sd7)^(-5'sd13))));
  localparam [4:0] p1 = {((-(+((4'd13)===(-3'sd0))))>(-((3'd4)?(-3'sd3):(2'sd1))))};
  localparam [5:0] p2 = ((~|(((-4'sd4)?(-5'sd13):(2'sd1))^((4'd11)^~(2'sd1))))?((~|(2'd2))|((-5'sd11)?(3'd6):(2'sd0))):(((-3'sd0)?(4'd6):(3'sd2))*((2'd2)+(5'd4))));
  localparam signed [3:0] p3 = {(!(|(-{(3'sd3),(2'sd0),(4'sd0)}))),{(&(4'd15)),{3{(2'd2)}},(+(5'd20))}};
  localparam signed [4:0] p4 = ((~^{2{(3'd4)}})<<{4{(4'd12)}});
  localparam signed [5:0] p5 = {1{{4{((4'sd3)?(3'd6):(3'd6))}}}};
  localparam [3:0] p6 = {3{{2{(3'd6)}}}};
  localparam [4:0] p7 = (3'd1);
  localparam [5:0] p8 = (~((^{4{(4'sd6)}})&{2{(-2'sd0)}}));
  localparam signed [3:0] p9 = (-{(~{(4'd5),(-4'sd7),(-3'sd3)}),{2{(4'd3)}},(-{2{(5'd3)}})});
  localparam signed [4:0] p10 = (~&((+(5'd26))*(~|(3'd0))));
  localparam signed [5:0] p11 = (5'd2 * (3'd0));
  localparam [3:0] p12 = (&(~&{4{(-3'sd1)}}));
  localparam [4:0] p13 = {1{((5'd28)?(4'd8):(-4'sd4))}};
  localparam [5:0] p14 = (~{(-(+({(3'sd2),(3'd6),(-5'sd6)}==(~|((5'd4)-(3'd0))))))});
  localparam signed [3:0] p15 = ((5'sd4)+(-3'sd1));
  localparam signed [4:0] p16 = {{((4'sd6)&&(4'd4)),(~&(4'd12))},(~|(~^(+{(2'd2)}))),(5'd2 * {4{(2'd3)}})};
  localparam signed [5:0] p17 = (((-3'sd1)!==(5'd18))?((-4'sd1)?(-5'sd6):(4'sd6)):((4'sd3)!=(2'sd1)));

  assign y0 = $signed((+p17));
  assign y1 = (-5'sd7);
  assign y2 = (~^{((4'd2 * p14)?(b2?b3:b5):$signed(p10)),(3'd6)});
  assign y3 = {((|({p13,p17,p6}<={4{b4}}))|(6'd2 * (p14<<a2)))};
  assign y4 = ({b4}&(~a2));
  assign y5 = (~|(+(-p4)));
  assign y6 = (~&(~&(!{2{((p1?p2:a5)?(p16?p13:p9):(p16?p11:p9))}})));
  assign y7 = (!(((|(~b4))*(a3>p4))&&((b5&b2)|(a4<<<a0))));
  assign y8 = {4{p14}};
  assign y9 = (2'd1);
  assign y10 = ((p7>=b5)||(b0>>>p2));
  assign y11 = (5'd1);
  assign y12 = $unsigned($unsigned(($unsigned((p10)))));
  assign y13 = ((&(p2^p0))||((|a1)||(~p13)));
  assign y14 = (((p16?p0:p3)/p17)?((p1<=p14)*(p1?p11:p4)):((p5>>>p16)+(p3?p1:p9)));
  assign y15 = (-(&($signed((^(~(p13>>>a0))))|(~&(|(!((a5))))))));
  assign y16 = {4{b2}};
  assign y17 = (5'd3);
endmodule
