module expression_00156(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'sd2)?((5'd15)>=(5'd21)):((4'd1)===(4'sd3)))>>({4{(2'sd0)}}-{4{(4'd2)}}));
  localparam [4:0] p1 = (!((4'd2 * ((2'd0)>>>(4'd11)))>>(3'd5)));
  localparam [5:0] p2 = (~^({4{(3'd6)}}?((-4'sd5)||(2'd2)):((-5'sd5)?(4'd6):(5'd4))));
  localparam signed [3:0] p3 = (+(~&{4{((3'd5)?(-2'sd0):(2'd1))}}));
  localparam signed [4:0] p4 = ({4{(4'sd5)}}===((3'd2)<(-3'sd2)));
  localparam signed [5:0] p5 = {{3{(~&((4'sd2)?(-2'sd0):(4'd12)))}}};
  localparam [3:0] p6 = (5'd2 * ((4'd2)===(4'd8)));
  localparam [4:0] p7 = (~(&(~&((-5'sd11)?(((-4'sd5)?(-3'sd0):(3'd2))==(&(5'd21))):(~&((2'd1)?(5'd6):(2'd2)))))));
  localparam [5:0] p8 = ((~&((5'd5)?(-2'sd1):(2'sd0)))?(((5'd23)?(-5'sd4):(3'd6))|((2'd0)?(3'd3):(4'sd4))):((~|(5'd7))===((5'sd9)*(5'd17))));
  localparam signed [3:0] p9 = (-2'sd0);
  localparam signed [4:0] p10 = ((-5'sd6)-(2'sd0));
  localparam signed [5:0] p11 = ((2'd1)>=(5'sd14));
  localparam [3:0] p12 = ({4{(3'd2)}}?{(5'sd8),(4'd12),(-3'sd3)}:((5'd19)<<(2'd3)));
  localparam [4:0] p13 = (((2'sd1)>>>(-5'sd14))>>>((2'd1)^~(-2'sd1)));
  localparam [5:0] p14 = (-(!(~^(2'd2))));
  localparam signed [3:0] p15 = ({((5'd6)+(-3'sd3)),((-3'sd3)===(-5'sd0)),((5'd19)<(3'sd0))}^~({(5'd22),(2'sd0)}===((-2'sd0)&&(5'd4))));
  localparam signed [4:0] p16 = {3{((-(4'd1))||((4'd5)^(3'd4)))}};
  localparam signed [5:0] p17 = ((3'd5)?((4'd12)+(-4'sd4)):((-2'sd0)?(3'sd3):(2'd1)));

  assign y0 = {(a4>a0),{3{a5}}};
  assign y1 = ((b4!==b0)>{b1,a3});
  assign y2 = (+(^(~|(~a5))));
  assign y3 = ((+{(!$signed((~^{p10,a2,a4}))),((~|(b0))|(a1+a2)),({(~|a1),{p17},(4'd2 * a1)})}));
  assign y4 = $unsigned((^(|(!{3{((p10^b3))}}))));
  assign y5 = $signed(((~(((!p6)>>(a2))>($unsigned(p3)>>{a4})))+(((a3&a2)===(b2===b3))<={(&a2),(~^b0)})));
  assign y6 = ((b2^b4));
  assign y7 = $signed($unsigned({$signed({p14,a3,b5}),(b5+p17),$signed($signed(a1))}));
  assign y8 = (((-a4)!=(b3?a4:p6))?(a4?p11:a4):(-(a1?b3:a0)));
  assign y9 = (|(-2'sd1));
  assign y10 = (b5?a4:a1);
  assign y11 = {(~(-{3{{p12,a1}}})),((~^{b0,p15})|{(p0^~a1)})};
  assign y12 = {2{(~^({2{(b1&&a1)}}==(~^(a4-a3))))}};
  assign y13 = (((p4!=p7)?(p17?p17:p12):(~p17))>=(-{(b5|p16),(p17?p1:p0)}));
  assign y14 = ((b4%b0)?$unsigned(p2):(p11+a3));
  assign y15 = (((-5'sd8)<<<((~^b1)<<<(a4&&b2)))>(4'd0));
  assign y16 = $unsigned(({3{{3{a4}}}}!==$unsigned(({2{b5}}?(b1-a2):(b3<<<a0)))));
  assign y17 = (~&{3{(-{3{a2}})}});
endmodule
