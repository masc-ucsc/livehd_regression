module expression_00698(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({((3'd7)>>>(2'd1)),((4'd5)!==(-2'sd0)),((4'sd6)^(3'd5))}&({(4'sd3),(3'sd2)}||((4'd7)-(-5'sd4))));
  localparam [4:0] p1 = ((&(4'sd7))===(^(-4'sd4)));
  localparam [5:0] p2 = (~(-{((-4'sd3)?(5'd15):(3'd6)),((2'sd0)?(2'd0):(-5'sd14))}));
  localparam signed [3:0] p3 = (((5'sd5)?(2'd0):(2'd0))?((4'd15)?(5'd6):(2'd3)):((2'd3)?(2'd1):(-2'sd0)));
  localparam signed [4:0] p4 = {2{{4{(-3'sd2)}}}};
  localparam signed [5:0] p5 = {(3'd0),(-4'sd2)};
  localparam [3:0] p6 = (4'd2 * (~^((4'd13)^(4'd0))));
  localparam [4:0] p7 = ({(3'd6)}|({(-3'sd2),(3'sd3)}<<{(3'sd0)}));
  localparam [5:0] p8 = (~^(&((~|{(4'd0)})^{((5'd26)<<(2'd3))})));
  localparam signed [3:0] p9 = (~((!(3'sd3))%(5'sd15)));
  localparam signed [4:0] p10 = (((-2'sd1)&(3'sd2))?((2'sd0)?(3'd4):(-4'sd3)):{(5'd10)});
  localparam signed [5:0] p11 = {3{{2{((2'd1)>=(2'd3))}}}};
  localparam [3:0] p12 = ({4{(2'd0)}}===((4'd12)?(2'd0):(-5'sd13)));
  localparam [4:0] p13 = (3'sd3);
  localparam [5:0] p14 = ((3'd3)*(-3'sd3));
  localparam signed [3:0] p15 = (~|(^{3{(^{4{(5'sd10)}})}}));
  localparam signed [4:0] p16 = (5'sd13);
  localparam signed [5:0] p17 = (^{1{(~(((3'd1)?(2'd0):(2'sd0))!==((-3'sd2)?(2'd1):(2'd3))))}});

  assign y0 = (((b2+p3)>>>{b3,a4,a5})>=({a4,p8}||{a1,b4}));
  assign y1 = ((~&p7)>=(p10<b4));
  assign y2 = ((-(p1<<<p11))!=(~(b0-p13)));
  assign y3 = ($signed(((a5?a1:b3)-(p3?b0:b0)))>=$unsigned(($signed((b3))||{3{b0}})));
  assign y4 = {1{((a5>>>b4)===(!{3{b4}}))}};
  assign y5 = {((~(~|a1))?{(2'd3)}:{b5,p10,b2}),((b0^b1)?(-{p3,b1}):(-{a5}))};
  assign y6 = {({1{(-5'sd11)}}!==(2'sd1)),(!((&p8)<<{2{p1}})),((~^p15)?(|p16):(p2?p1:p14))};
  assign y7 = {{1{{1{{4{{{2{a1}}}}}}}}}};
  assign y8 = {4{(-(4'sd1))}};
  assign y9 = (($signed($signed((p12>a3)))^~((p16>p8)||$signed(p12)))^~((((p6<<p16)|(a5===b0))^$unsigned($unsigned((p6==p12))))));
  assign y10 = $signed((((((5'sd1))|(2'd0))^{{p10,a2,b4},$signed((a1|a0))})));
  assign y11 = (!p17);
  assign y12 = ((3'sd3)<({p4,a5}-(&b3)));
  assign y13 = (({(|{(|a4)})}&&(~|{(a5-b3),{b3,a4,p0}}))>>>{(~({{a4,b4},(~|b2)}!==(-{(a1||a5)})))});
  assign y14 = ((a5?a2:a1)?(a1?b3:b4):(&(a2?b3:a3)));
  assign y15 = (|{(!(~^(p17?p14:p9))),{(p0?p16:p1),(p16?b2:p14)}});
  assign y16 = ({4{{2{p6}}}}==(({4{p16}}&&(p9+p6))>>>((p16>=p0)>>(a5!==b1))));
  assign y17 = {1{(~&((|{{1{{a1,a2,b3}}},(a5?b1:a3)})!==((&(~b1))?{(!a2)}:(b1!=a4))))}};
endmodule
