module expression_00071(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{((2'd2)?(2'd3):(4'd8))},(2'd0)};
  localparam [4:0] p1 = ((-4'sd4)?(5'd5):(2'd3));
  localparam [5:0] p2 = (((5'd6)>>(2'd3))<<((5'sd7)!=(3'sd0)));
  localparam signed [3:0] p3 = ({(|(3'd7)),{1{(2'd2)}},(+(-2'sd1))}-{((-5'sd14)!=(-5'sd10)),{4{(4'd10)}},{(5'd22)}});
  localparam signed [4:0] p4 = (4'sd6);
  localparam signed [5:0] p5 = (|(~|(+(&(!(~(&(~&(~^(&(2'sd1)))))))))));
  localparam [3:0] p6 = (((((4'sd5)?(2'sd1):(-4'sd2))<<{2{(-3'sd0)}})&((2'sd1)?(-4'sd7):(3'd6)))&(~^((5'd2 * (5'd5))||((2'd3)^~(4'sd3)))));
  localparam [4:0] p7 = (((2'd2)==(3'd2))*(^(4'd8)));
  localparam [5:0] p8 = {4{{(5'd4),(4'd15),(3'sd0)}}};
  localparam signed [3:0] p9 = (4'sd3);
  localparam signed [4:0] p10 = {{(2'sd1),(4'sd6),(-5'sd7)},((5'd19)&(4'd0)),(-5'sd8)};
  localparam signed [5:0] p11 = ({2{((3'sd1)>>(3'd6))}}||{4{((3'd1)!=(-2'sd1))}});
  localparam [3:0] p12 = {1{((-(-4'sd7))+(-(-4'sd4)))}};
  localparam [4:0] p13 = (5'sd5);
  localparam [5:0] p14 = {3{(((4'd9)?(4'd14):(5'd23))<{2{(2'd3)}})}};
  localparam signed [3:0] p15 = (((2'd3)?(2'd2):(5'd5))?{(-2'sd1),(5'd21)}:((-2'sd0)==(2'sd1)));
  localparam signed [4:0] p16 = ((2'd3)?(5'sd2):(-4'sd6));
  localparam signed [5:0] p17 = ((|((2'd2)<<(-4'sd6)))/(2'd2));

  assign y0 = (((b1!=p7)==(b3>>a2))>>>((b2|b3)&&{b0,a0,a0}));
  assign y1 = ((((a1<=p17))>={(~^a4)})<<<({b3,b2}<<<(p14+b5)));
  assign y2 = (((a0)==={3{a2}})|{a3,a5,a0});
  assign y3 = $unsigned(($signed(a4)?(p6?p8:a4):(p17?a2:p5)));
  assign y4 = $unsigned({{(-2'sd0),(b1>>>b1)}});
  assign y5 = (4'd15);
  assign y6 = {1{({a0,b4}?{a5,b5,a4}:{3{a5}})}};
  assign y7 = (((~^p9)&&{b5})?{1{{4{p17}}}}:{($unsigned(p4)|{b1,a4})});
  assign y8 = {2{{1{(5'd29)}}}};
  assign y9 = (((a3?a0:b0)&&(a3<<b0))<<((b3!==a0)==(+(a0>>>b1))));
  assign y10 = (~^((2'sd1)<=(2'sd1)));
  assign y11 = (5'd7);
  assign y12 = (2'd1);
  assign y13 = (|(a3+a0));
  assign y14 = {(b1?a1:a4),{(~|b4)},(-(p16?b2:p4))};
  assign y15 = (5'sd3);
  assign y16 = (-(-5'sd1));
  assign y17 = $signed($unsigned(((({3{p15}}>>>(p13))?(5'd13):{3{p9}}))));
endmodule
