module expression_00811(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd3);
  localparam [4:0] p1 = (+((4'd2 * (4'd0))?(~&(~|(2'sd0))):{(5'd7),(-2'sd1),(-2'sd1)}));
  localparam [5:0] p2 = (^(-5'sd9));
  localparam signed [3:0] p3 = (((-2'sd1)?(-4'sd5):(-4'sd7))/(-2'sd1));
  localparam signed [4:0] p4 = ((4'sd4)?(5'sd13):(-4'sd4));
  localparam signed [5:0] p5 = ((((2'd3)?(5'd18):(2'd3))?((3'sd1)?(4'd8):(5'd11)):((5'd6)>>>(5'd10)))|(((3'd6)?(3'd7):(-5'sd3))==(((4'd1)-(3'd0))>{(4'd12),(-2'sd1),(4'd8)})));
  localparam [3:0] p6 = (-3'sd0);
  localparam [4:0] p7 = (-{1{({3{((-3'sd0)<(3'd6))}}<{3{((3'sd1)<(3'sd3))}})}});
  localparam [5:0] p8 = (((2'sd1)?(5'd22):(4'd4))|((2'd2)>>(-2'sd0)));
  localparam signed [3:0] p9 = ((((4'sd3)==(5'd25))===((-4'sd2)&(3'sd3)))^(((5'sd1)|(2'sd1))>=((5'sd13)!=(-4'sd0))));
  localparam signed [4:0] p10 = ((~|((3'd3)!=(5'd8)))^~(!(^((3'd4)%(4'd0)))));
  localparam signed [5:0] p11 = (((4'sd4)>(-5'sd0))!=((-2'sd0)<<<(-4'sd6)));
  localparam [3:0] p12 = (^(5'd18));
  localparam [4:0] p13 = (((5'd2 * (2'd2))>{(4'sd3),(5'd19),(4'sd2)})>{{(2'sd1)},{(2'd2),(3'd1),(-3'sd3)}});
  localparam [5:0] p14 = ({3{(2'sd0)}}+(-(3'd5)));
  localparam signed [3:0] p15 = (^((-4'sd4)?((2'sd0)?(3'd6):(-4'sd7)):((2'sd1)?(4'sd1):(-3'sd1))));
  localparam signed [4:0] p16 = ((&(5'd11))?((3'd3)?(5'd14):(2'sd0)):{2{(2'd1)}});
  localparam signed [5:0] p17 = (((3'd7)?(4'd2):(4'sd2))%(3'sd3));

  assign y0 = (~&(~^$signed((~^(~^(~&$unsigned($signed(a4))))))));
  assign y1 = ($unsigned((-5'sd10))==(^((2'd2)>=((b4+a3)))));
  assign y2 = (4'd11);
  assign y3 = ((3'd3)?(-5'sd9):(p7?a0:a2));
  assign y4 = ((!(!(~(|(~(&(-(p9<<<a2))))))))>(+((!(6'd2 * a0))!==(~(!(~&a5))))));
  assign y5 = {a4,p11,a1};
  assign y6 = {1{{1{((($unsigned((a5===b0))|(b3?p1:a3)))+((b2?b4:p1)&&(a0>b5)))}}}};
  assign y7 = ((&{{p10},(p1?p11:p5)})>((6'd2 * p1)|{3{a3}}));
  assign y8 = ((((b0>a2)!==(a5<<<b5))>=(!(^(b1<=a3))))>>((p8?a3:p6)>>((b0?p12:a1)^~(~^b4))));
  assign y9 = {3{b5}};
  assign y10 = (((a2|b2)!=(6'd2 * a1))===((a5-b1)==={3{b2}}));
  assign y11 = (|{2{{2{a5}}}});
  assign y12 = ({a2}^(a2&p17));
  assign y13 = (5'd28);
  assign y14 = (-(~&(4'd4)));
  assign y15 = ({(a1?p2:b5),{p15},(-3'sd0)}?{((b3?b2:a3)?(b2?b5:p13):(b2?a3:p16))}:{(a1?a0:p4),{b4,b4,a0},{b3,b0}});
  assign y16 = ($unsigned($unsigned($signed(($unsigned(a3)?(b4^b0):(a0?p14:a5))))));
  assign y17 = ({2{p10}}<(~&a0));
endmodule
