module expression_00775(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&((-3'sd3)?(5'd8):(4'd9)));
  localparam [4:0] p1 = ({2{(3'd1)}}?((4'd10)>>(-3'sd0)):((4'd11)?(3'd6):(-5'sd6)));
  localparam [5:0] p2 = ((3'sd3)^(4'd14));
  localparam signed [3:0] p3 = {1{(2'sd1)}};
  localparam signed [4:0] p4 = {{2{(5'd22)}},{(2'd1),(5'd23),(4'd8)}};
  localparam signed [5:0] p5 = ((((4'd11)&(2'd0))>>>((-5'sd2)?(2'sd0):(4'd2)))&&{(((4'd9)?(4'sd7):(5'sd2))+{(3'd7),(4'd12),(3'd2)})});
  localparam [3:0] p6 = {3{(!({(2'sd0),(2'd0),(-3'sd0)}+{2{(5'sd15)}}))}};
  localparam [4:0] p7 = ((3'd0)?(|(2'sd1)):({1{(-2'sd1)}}?((-4'sd0)?(2'd3):(2'sd1)):(5'd12)));
  localparam [5:0] p8 = {((2'd1)<<(-5'sd12))};
  localparam signed [3:0] p9 = ((-2'sd1)^~((3'd3)!==(-4'sd3)));
  localparam signed [4:0] p10 = (&(((4'd7)>=(2'd2))^(^{(-4'sd3),(2'd3),(4'd4)})));
  localparam signed [5:0] p11 = (&((!(-(-2'sd1)))?(-((2'd3)?(5'sd4):(5'd19))):(~^(~(5'd10)))));
  localparam [3:0] p12 = ((((4'd2)?(5'sd2):(4'd12))?((-5'sd7)^~(5'd23)):((4'sd6)?(2'd0):(-4'sd1)))&&(((4'sd2)<<<(2'd0))!=((-3'sd0)?(4'd3):(4'sd4))));
  localparam [4:0] p13 = (~^(^(+((-2'sd1)>=(3'd0)))));
  localparam [5:0] p14 = (~((((3'd3)&(2'sd1))<={(|(4'sd3))})!==(~^(+((+(3'd4))?((5'sd11)?(2'd1):(5'sd10)):(+(2'd2)))))));
  localparam signed [3:0] p15 = ({((-4'sd2)?(4'sd3):(-3'sd1)),((2'd3)?(4'd4):(3'd7))}===(~|((-4'sd3)?(3'd1):(-4'sd1))));
  localparam signed [4:0] p16 = ((~^((5'd26)&(2'd2)))>>>(~|(~(2'd0))));
  localparam signed [5:0] p17 = ((-4'sd7)>>>(+((2'd0)?((-5'sd0)?(2'sd1):(2'd0)):(-(4'd6)))));

  assign y0 = ((~|p12)+(-4'sd6));
  assign y1 = ({3{a2}}?(!p17):(p16?a4:a2));
  assign y2 = {(-2'sd1),(-4'sd1),(5'd0)};
  assign y3 = (((~^b1)>>>{4{a5}})?({4{a5}}?(a1+b1):(a1?a3:a2)):((a0<b2)?{1{b5}}:{1{a3}}));
  assign y4 = (^{4{{p15,a5,p2}}});
  assign y5 = ({(a4!==b5),{p10,p12}}&($signed(b3)&$signed(p7)));
  assign y6 = ((~p12)!=(-2'sd1));
  assign y7 = ((((b2>>>p0))>=(-3'sd1))||((a1<=p14)?(a2<=p4):(p12?p11:p17)));
  assign y8 = (^p4);
  assign y9 = (5'd2 * (-(p6<<p12)));
  assign y10 = ($signed(((p6||p0)>$unsigned(p11)))>>>((p4)==(p16==p14)));
  assign y11 = {b4,b0};
  assign y12 = {2{(p11?a4:b3)}};
  assign y13 = {3{{2{b4}}}};
  assign y14 = ({3{(b4)}}<<<({1{(a2+a1)}}!=$signed($signed(b4))));
  assign y15 = (5'd2 * {1{(a0&&a2)}});
  assign y16 = (~|(3'd5));
  assign y17 = {$signed($unsigned({3{(p1)}})),{{p13,b4,p5},{p8,b0,a3}},(~(({b4}?(!b4):(p15?p13:a3))))};
endmodule
