module expression_00017(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd0)>=(2'd0))^~(^((4'sd4)?(-5'sd12):(2'sd0))));
  localparam [4:0] p1 = ({1{(-5'sd0)}}<<{1{({1{(-2'sd1)}}>>>((4'd12)|(3'd0)))}});
  localparam [5:0] p2 = ((-(4'd2 * (-(2'd3))))>>>(((4'd4)&(2'd2))&&((-5'sd8)*(4'd14))));
  localparam signed [3:0] p3 = ((5'd2 * (3'd0))^~(6'd2 * (2'd3)));
  localparam signed [4:0] p4 = (((3'd0)<<<(-5'sd5))?((4'd0)>>(2'd3)):((5'd18)?(5'd0):(4'd4)));
  localparam signed [5:0] p5 = (-(!((~(-3'sd0))<((2'd2)&&(-4'sd7)))));
  localparam [3:0] p6 = (({(2'sd0),(5'd8),(5'sd11)}<<{((-2'sd1)&(-2'sd1))})&(4'd3));
  localparam [4:0] p7 = (~|((-(5'd21))?((4'd2)>>>(2'd1)):((2'd3)<<<(5'sd0))));
  localparam [5:0] p8 = (-{3{(4'd4)}});
  localparam signed [3:0] p9 = {1{((2'sd0)>>>(^(-5'sd7)))}};
  localparam signed [4:0] p10 = (~^(~(~{(3'sd1)})));
  localparam signed [5:0] p11 = (-5'sd0);
  localparam [3:0] p12 = (^((4'sd7)^(2'd2)));
  localparam [4:0] p13 = ({4{(5'd6)}}?{1{(2'sd1)}}:{3{(-2'sd1)}});
  localparam [5:0] p14 = {(&((-4'sd1)?(4'd5):(3'd5))),((5'd11)?(-4'sd5):(-4'sd4)),((2'd1)?(2'd3):(-3'sd0))};
  localparam signed [3:0] p15 = (^(~(-4'sd5)));
  localparam signed [4:0] p16 = ({4{(-3'sd2)}}|((4'sd6)||(-2'sd1)));
  localparam signed [5:0] p17 = ({1{(3'd3)}}?((4'd10)^~(3'd7)):((-4'sd7)>>(-3'sd2)));

  assign y0 = ({(&p1),(^p16),(&p14)}>(^(~|((p6&p7)?(p7?p1:p10):(|p0)))));
  assign y1 = ((({1{p1}}-(4'd14))>=({1{b1}}+(2'sd1)))^~((a5^~p17)?(a3|p14):(b5<=a2)));
  assign y2 = ((((a0!==b3)+(6'd2 * p8))^(!{2{a4}}))<{1{({3{p8}}|(|{3{p0}}))}});
  assign y3 = (~(-{2{p2}}));
  assign y4 = {2{({4{p5}}&&(p15||p6))}};
  assign y5 = {1{((3'd2)?(-2'sd1):{(p6?p1:p15),(2'd0),(p16?p15:p3)})}};
  assign y6 = (+{(|(+{p0,p3})),{{2{p14}},{p9,p7}},{p4,b4,p1}});
  assign y7 = {(^{2{p14}})};
  assign y8 = (~&b2);
  assign y9 = ({4{$unsigned(a1)}}!==((b2?b2:b5)?(a0?a4:b3):(a0!==a0)));
  assign y10 = $signed({({p7,a1}>>>$unsigned(p16)),$signed(((p13>b1)&&(2'sd0)))});
  assign y11 = (&{4{{4{b3}}}});
  assign y12 = $unsigned($unsigned(((~^(-p0))==(!$signed(b1)))));
  assign y13 = ((-3'sd2)<{4{b4}});
  assign y14 = ((-(a3?b0:p11))?{p9,p6,p7}:{a1,p9});
  assign y15 = ({3{(p14==b4)}}<<<(~|{3{(^a5)}}));
  assign y16 = ({1{((a0!=b3)<<<{1{b0}})}}>((p15>>b0)&{2{p3}}));
  assign y17 = (~($unsigned((~^$unsigned((!(~&$unsigned(((-(-$signed((&(p1))))))))))))));
endmodule
