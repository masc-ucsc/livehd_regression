module expression_00205(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(((3'sd3)<(2'sd1))!==(4'sd6))}};
  localparam [4:0] p1 = (((-5'sd11)?(3'd6):(2'sd1))?((5'sd8)?(4'sd3):(5'd15)):((-2'sd0)?(5'd7):(4'd8)));
  localparam [5:0] p2 = (((5'd6)>>(2'd1))>>((2'd1)/(3'sd1)));
  localparam signed [3:0] p3 = ((5'd9)||(-5'sd11));
  localparam signed [4:0] p4 = (~^(~(&(((5'd9)===(3'sd2))!={{(5'sd5)}}))));
  localparam signed [5:0] p5 = ((~|{{(3'sd2)}})^({{(2'd3),(4'sd7),(-2'sd1)},((-3'sd1)<<<(5'sd10))}<<{((2'sd0)+(3'd1)),{(3'd4),(4'sd4),(3'sd1)}}));
  localparam [3:0] p6 = {2{{3{(3'd0)}}}};
  localparam [4:0] p7 = {4{{4{(2'sd0)}}}};
  localparam [5:0] p8 = (2'd3);
  localparam signed [3:0] p9 = {3{((-2'sd0)?(-5'sd2):(5'd11))}};
  localparam signed [4:0] p10 = ({{{3{(-4'sd5)}}},(~|((-5'sd1)<<(2'd3)))}<<<{2{(-((2'd0)-(4'd2)))}});
  localparam signed [5:0] p11 = {(2'd2),{2{((5'd1)>=(2'sd1))}},{(2'd3),(2'd3),(3'd4)}};
  localparam [3:0] p12 = ({3{(~{1{(4'sd2)}})}}>>>(-2'sd0));
  localparam [4:0] p13 = (((-4'sd0)===(4'sd5))?((3'sd0)+(4'sd5)):((-4'sd1)?(4'sd6):(3'd6)));
  localparam [5:0] p14 = (~&{3{(((-5'sd2)&(2'd0))<=(~|(5'd10)))}});
  localparam signed [3:0] p15 = (^{1{(!{3{(2'd2)}})}});
  localparam signed [4:0] p16 = {{{1{(-((5'd8)&&(5'd6)))}},(4'd2 * ((4'd10)-(2'd3)))}};
  localparam signed [5:0] p17 = (((((5'sd8)*(-3'sd3))==((2'sd1)>(4'd3)))+((5'sd0)%(-2'sd1)))>((((5'd8)!==(4'd12))||((2'sd1)!=(4'sd0)))<<(((3'd0)|(-3'sd1))||((4'd7)<<(4'd4)))));

  assign y0 = ({3{$unsigned(b0)}}<<({4{p2}}!={4{a2}}));
  assign y1 = (2'd1);
  assign y2 = ((!p10)>>>(~&p17));
  assign y3 = (((-(^(+(~^b0)))))?(&(~&(&(!{3{p5}})))):($signed(p3)?(b2?p13:p17):(~&p13)));
  assign y4 = ((2'd2)?(^(~{3{p12}})):{2{(4'sd2)}});
  assign y5 = $signed({(5'd0)});
  assign y6 = (((~|p13)^~(p7%p10))-(~($unsigned(a0))));
  assign y7 = ($unsigned(p10)?(b2?a3:p15):(a5));
  assign y8 = ($unsigned((|(((p6?p10:p6))^((~&p10)==(a3-p16)))))<<(~&{((p6&a5)?$signed((~|a0)):(~^(a5?p0:p11)))}));
  assign y9 = (~|$unsigned((!{4{(+b4)}})));
  assign y10 = {(-2'sd0),(3'd3)};
  assign y11 = (4'd2 * $unsigned((|a5)));
  assign y12 = {3{(~^(^{3{p2}}))}};
  assign y13 = ({a1,a4,a0}===({b4}&{b5,b3,a4}));
  assign y14 = ((4'sd2)>=((p11-p15)&(p5?p3:b0)));
  assign y15 = {((!b1)||(p8?b5:b2)),{(4'd2 * (&a0))},((a1?b5:b2)?(b1?b1:a5):(b0!==a0))};
  assign y16 = ((5'd2 * p13)!=(4'sd4));
  assign y17 = ((~^{1{{3{(-a2)}}}})===(-({b1,a0,a0}|{(b3^b2)})));
endmodule
