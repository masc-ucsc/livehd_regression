module expression_00881(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd2);
  localparam [4:0] p1 = {({(5'd13)}|{(4'd5),(2'd3)})};
  localparam [5:0] p2 = ({(-5'sd10),(3'd2),(-3'sd2)}?(~&(4'sd3)):{(-4'sd5),(-4'sd4),(4'd5)});
  localparam signed [3:0] p3 = {4{((3'sd0)^~(-4'sd3))}};
  localparam signed [4:0] p4 = (-2'sd0);
  localparam signed [5:0] p5 = {{4{(4'sd1)}}};
  localparam [3:0] p6 = ((4'sd5)^~((4'd14)<(3'd6)));
  localparam [4:0] p7 = ((~&(~|(3'd1)))-((4'd6)||(3'd5)));
  localparam [5:0] p8 = ((-({(-3'sd3),(2'd0),(-4'sd2)}!=((4'd0)^~(4'd4))))>=(((2'd1)<=(3'd1))&&((-5'sd5)>(3'd2))));
  localparam signed [3:0] p9 = (~&(~|(^((^{1{(-4'sd0)}})?(!((-4'sd2)+(-4'sd3))):((4'd2)&&(-3'sd2))))));
  localparam signed [4:0] p10 = ((5'd13)?(-5'sd13):((4'd9)>(2'sd1)));
  localparam signed [5:0] p11 = ({2{(2'd3)}}||((-4'sd4)>=(5'd16)));
  localparam [3:0] p12 = ((((4'sd1)^~(4'd6))<<<{(4'd14)})?(((4'd11)^(4'sd5))+((4'sd5)-(2'd0))):(~^{(-5'sd8),(-5'sd0),(-4'sd0)}));
  localparam [4:0] p13 = (-5'sd13);
  localparam [5:0] p14 = (~&(&{(5'd20),(3'sd2),(-3'sd1)}));
  localparam signed [3:0] p15 = (-(~|((3'sd2)^~(-5'sd11))));
  localparam signed [4:0] p16 = (^(~&(((^(5'd25))&((2'sd0)+(2'd0)))?((!(-3'sd0))||{(-3'sd3),(3'sd0)}):(-((5'd12)<<(3'd7))))));
  localparam signed [5:0] p17 = ((-5'sd2)?(2'd0):(4'sd2));

  assign y0 = {(4'sd6),((a1|b4)&&(b3!=p10)),$unsigned((~|(p9)))};
  assign y1 = {4{((!p1)?$signed(p17):$signed(p1))}};
  assign y2 = ((~|(b0<<a5))?(~(a2===a1)):{p16,b0,p13});
  assign y3 = ((2'd0)||(-(~(6'd2 * (^b0)))));
  assign y4 = ((+p0)?(p7):(b3&b4));
  assign y5 = (2'd1);
  assign y6 = (p6?p5:p14);
  assign y7 = (&(-2'sd0));
  assign y8 = {1{$unsigned(((-3'sd2)<(b5+p9)))}};
  assign y9 = ((p15||p3)%p0);
  assign y10 = (((a4|b4)?(b1?b2:b0):{3{b5}})===$signed((b5?a2:a5)));
  assign y11 = {1{(~&a1)}};
  assign y12 = $signed((5'd14));
  assign y13 = (((p16<<p3)||(p4>>p3))>>>((p6>p4)>(p7&&p3)));
  assign y14 = {{(a3),{p2,p17,p7}},$signed((p5|b0)),{(p4+b4)}};
  assign y15 = $signed($unsigned(p5));
  assign y16 = (b5?a2:b0);
  assign y17 = (($unsigned($signed((a3>p14)))>$unsigned({p8,b0,b1}))>>$unsigned(($signed({a2,b2})||($unsigned($signed(a2))))));
endmodule
