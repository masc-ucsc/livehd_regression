module expression_00316(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(&((3'd5)>>(5'd16)))}};
  localparam [4:0] p1 = (2'd3);
  localparam [5:0] p2 = ((3'sd0)^(2'd1));
  localparam signed [3:0] p3 = (~^((!(~^({2{(-3'sd3)}}?((-3'sd0)?(2'd0):(-2'sd0)):(+(-5'sd3)))))^(((5'd10)!=(-5'sd4))<((5'd17)>(3'd4)))));
  localparam signed [4:0] p4 = ((-((~&((-3'sd0)>>(5'sd10)))<<<((4'sd4)<(-5'sd0))))>>>(((-3'sd0)||(5'd15))?((2'sd0)>=(-3'sd2)):((-3'sd0)!==(4'd0))));
  localparam signed [5:0] p5 = {4{((-5'sd13)>(-2'sd0))}};
  localparam [3:0] p6 = (~&((4'sd3)||(2'sd1)));
  localparam [4:0] p7 = (~^{2{(4'sd6)}});
  localparam [5:0] p8 = ((5'd2 * (2'd2))*(|(5'd7)));
  localparam signed [3:0] p9 = ((4'd10)<<<(-5'sd6));
  localparam signed [4:0] p10 = (~|{{{(5'sd10),(3'sd3)},{4{(2'd0)}},{1{(-4'sd2)}}},{{(2'd3),(3'd5),(4'd15)},((-5'sd4)>>>(3'd1)),(2'sd1)},(4'd1)});
  localparam signed [5:0] p11 = (!{(((-4'sd7)?(5'd6):(4'd8))&{4{(-3'sd1)}})});
  localparam [3:0] p12 = ((-3'sd3)<=((2'd3)==(-5'sd4)));
  localparam [4:0] p13 = (-{((5'd6)^(3'sd3)),(|(4'd5)),{4{(2'd0)}}});
  localparam [5:0] p14 = (~|((-4'sd4)&(3'sd0)));
  localparam signed [3:0] p15 = {3{((5'd28)?(4'sd5):(3'sd0))}};
  localparam signed [4:0] p16 = (|{3{(&(~(-2'sd1)))}});
  localparam signed [5:0] p17 = (~|(5'd6));

  assign y0 = {{b3,a3,a0},(a5|b5)};
  assign y1 = $signed(p1);
  assign y2 = (-((~^{$unsigned(b3),(p8?p5:p3)})?$unsigned((4'sd3)):((p16>p5)?$signed(p12):{p4,p0})));
  assign y3 = {{p4,p10},(b0?b5:b1),{$unsigned(b2)}};
  assign y4 = {4{(~|(a3^~b5))}};
  assign y5 = (2'd0);
  assign y6 = {{$unsigned(b5),{b5,b2,b3},(4'sd1)},(-2'sd1)};
  assign y7 = {1{({1{{1{(~^(^{2{p12}}))}}}}<(!(^(~&(&{1{(p11!=p8)}})))))}};
  assign y8 = ({3{a4}}?(&(+b4)):(p15<b4));
  assign y9 = (($unsigned({(~|(+$signed({b4,p3,p4})))})||(5'd2 * (p1-p14))));
  assign y10 = ((((p5&b1)<<<(b5+p9))|((b0>>>p0)%p1))&(((b2>=a5)!=(p15<=p17))+((p4%p3)^(p2<b3))));
  assign y11 = $signed((^(((~|(p8-p0))>>(!(p1>p12)))|((&(p8^~a2))<=(a3/p3)))));
  assign y12 = (5'sd7);
  assign y13 = (~|(~^((b4&&b2)<<<(^(~&a0)))));
  assign y14 = (!(((b4!==a3)!=(p10>=a0))&(^(~^$signed(p7)))));
  assign y15 = ({(p7?p17:p6)}?{(b0!==a4),(p7?p14:p13)}:((p17|p10)||(p16<=p14)));
  assign y16 = {(~&p8),(a3!==b1)};
  assign y17 = (~$unsigned((~|(~(({3{p3}}<<(~(b2||a3)))<<((&(~|(~|b1)))==((p11+p10)>={1{p8}})))))));
endmodule
