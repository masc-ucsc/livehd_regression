module expression_00460(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd27)<<<(-4'sd6));
  localparam [4:0] p1 = ((((5'sd1)!==(3'sd1))&&((2'd2)?(2'd0):(-5'sd6)))<(((2'd1)&&(-3'sd1))>>>((4'sd7)&(2'sd0))));
  localparam [5:0] p2 = ((((-4'sd7)<=(-2'sd1))>(!(+(2'd1))))>>>(|(&((!(2'sd1))>(+(-5'sd1))))));
  localparam signed [3:0] p3 = {1{(~|(~^((-2'sd0)>(2'd0))))}};
  localparam signed [4:0] p4 = ((2'd0)-(4'd3));
  localparam signed [5:0] p5 = {3{{3{{1{(2'sd1)}}}}}};
  localparam [3:0] p6 = ({2{(3'd5)}}<<<((5'sd12)==(2'd3)));
  localparam [4:0] p7 = ({(2'sd0)}=={{(4'sd7),(5'd14),(-2'sd1)},{(2'd3),(2'd3)}});
  localparam [5:0] p8 = (5'sd15);
  localparam signed [3:0] p9 = ({3{(3'sd0)}}?(((3'd3)!=(2'sd1))?(&(4'd14)):{2{(2'd2)}}):({4{(2'sd0)}}?(-5'sd0):(~&(2'd3))));
  localparam signed [4:0] p10 = {4{(-4'sd4)}};
  localparam signed [5:0] p11 = ({(2'd3)}<=((5'd0)&&(-4'sd6)));
  localparam [3:0] p12 = (((5'd15)+(-4'sd5))*(-2'sd0));
  localparam [4:0] p13 = {(-2'sd0)};
  localparam [5:0] p14 = (4'sd0);
  localparam signed [3:0] p15 = (5'd1);
  localparam signed [4:0] p16 = (6'd2 * ((2'd3)<<<(3'd2)));
  localparam signed [5:0] p17 = {{((-3'sd3)>>>(5'd2)),((3'd7)===(3'd6)),(~&(-4'sd6))},(&{(~^((5'sd7)===(5'sd3)))})};

  assign y0 = (-5'sd12);
  assign y1 = (~&{3{{2{p4}}}});
  assign y2 = ({1{((|(a2-a5))>($unsigned(b2)!==(~|b0)))}}||($unsigned((a0^b4))^~((~&b5)|(b0))));
  assign y3 = (5'sd14);
  assign y4 = {($unsigned(p8)==(b0?p10:p14)),((b4>>>a1)-{b0}),(p1?a0:p9)};
  assign y5 = ((b5===b5)!=(p17<<p8));
  assign y6 = ($signed((+{1{(-p14)}}))<<((!p12)^~{p3}));
  assign y7 = (&{1{{3{(2'sd1)}}}});
  assign y8 = {2{{1{{(p4?p0:p7)}}}}};
  assign y9 = (((b0|a0)<<(b4>>>a3))^((b0>>a4)-(b0/b1)));
  assign y10 = (((+p8)>>(5'd24))-(5'sd10));
  assign y11 = ((+((^(p3+p2))!=(~&{1{p17}})))<{2{{2{(&p8)}}}});
  assign y12 = (^(~^{(p16?p7:p15),(~&a4),(-p17)}));
  assign y13 = {(a4!==a5),(~|p7)};
  assign y14 = (~^{2{(~|(^p3))}});
  assign y15 = (p8==a0);
  assign y16 = $signed((-5'sd1));
  assign y17 = $unsigned({2{b3}});
endmodule
