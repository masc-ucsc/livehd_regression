module expression_00653(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd3)?(-2'sd1):(3'd2));
  localparam [4:0] p1 = {(&{{{(3'd6)},{(5'd12)},(|(4'd5))},{(^(2'd2)),((5'sd2)===(5'sd13)),((-2'sd0)>>>(2'sd0))}})};
  localparam [5:0] p2 = ((((3'd3)==(5'd13))>((3'sd1)^~(5'd30)))!=(((3'd0)^(-3'sd1))&((2'sd0)<=(-4'sd2))));
  localparam signed [3:0] p3 = (-(!((5'd11)?(5'd1):(5'sd7))));
  localparam signed [4:0] p4 = (+{(~^(|{3{{(4'sd5),(5'd1)}}}))});
  localparam signed [5:0] p5 = {{(2'd1),(3'd1)},{(5'd24),(3'sd0)},((5'd6)===(5'd20))};
  localparam [3:0] p6 = {(((2'sd0)|(2'd2))&((2'sd1)>=(2'd0))),(~&(4'd2 * (3'd1)))};
  localparam [4:0] p7 = (+(3'd7));
  localparam [5:0] p8 = (((2'sd0)<=(4'd12))>>((-3'sd3)>(-2'sd1)));
  localparam signed [3:0] p9 = (((5'sd15)|(^(5'd2 * (3'd6))))^~(-(~(4'sd0))));
  localparam signed [4:0] p10 = ((5'd14)?(3'd6):(((-5'sd14)^(5'd29))>(4'd15)));
  localparam signed [5:0] p11 = (^(((4'sd6)>>((4'd5)&&(2'd0)))^(-3'sd2)));
  localparam [3:0] p12 = (((2'd1)*(3'sd1))<(|((5'd5)<(2'sd0))));
  localparam [4:0] p13 = (~((-2'sd1)?(5'sd3):(5'd25)));
  localparam [5:0] p14 = ((3'sd0)!==(((4'd0)<<(2'd1))<<<((-3'sd2)+(4'd2))));
  localparam signed [3:0] p15 = {1{{4{(2'd2)}}}};
  localparam signed [4:0] p16 = ((-4'sd5)==(2'sd0));
  localparam signed [5:0] p17 = {(-2'sd0),(-5'sd3),(4'sd2)};

  assign y0 = $unsigned({3{$signed((~(p11&&p11)))}});
  assign y1 = (+(~^(~^(~&(~^(!(~&(!(~^(|(|(~|(&(&(~|(!(!p13)))))))))))))))));
  assign y2 = {({(p15<=p11)}-{(p16<<p15)}),{(a1<p0),(p13+p15),(p8<=b5)}};
  assign y3 = ($unsigned(({3{a4}}>>(p8)))?((p11&a5)?(p10?a5:p6):(p5<=p5)):({3{p8}}||(b0<=a3)));
  assign y4 = (-((4'd2 * (b2&&b0))<((p14?a2:p15)?(a0===a4):((a0===a1)))));
  assign y5 = {2{a3}};
  assign y6 = (((a5-p1)>>>(a4^~b1))<<{1{((a3>>p4)!={4{b0}})}});
  assign y7 = ({a5,a4,b2}?$unsigned((b4?a1:b4)):$unsigned((b0?a4:a2)));
  assign y8 = (~&((|(+(b0^p4)))>>>{{4{p9}},(&b0)}));
  assign y9 = ((2'sd1)>$unsigned((+$unsigned(b4))));
  assign y10 = ({(!{a4}),(~(&p15)),{b1,p12,a1}}>>{(^{$signed(b0)}),{(+p2),$unsigned(a3)}});
  assign y11 = {4{(b3<=a2)}};
  assign y12 = (p16?p11:p14);
  assign y13 = (~((((a0*p16)<<(-4'sd1))&&(((+b3))))<=$signed((+(((b3===b1))/p13)))));
  assign y14 = ((({p12,p3}>>{p15,p4})>=({p15}?{p17,p17}:(p4?p12:a0)))<<<(((5'd7)?(p11?p6:p12):{a0,a1,a3})<=((a1==p4)?(p10?p5:p2):(p16?p14:p2))));
  assign y15 = ($signed($signed((((a4||a1))===((a5==b4)^(b5&&b2)))))>$unsigned((((b3===a1)>=(a4))!=((a1<<p15)-(p0*b1)))));
  assign y16 = (((b5-b5)<<<{b5,b3,a1})<(^{b4,b4}));
  assign y17 = (+(!({p8,b4}?(-2'sd1):(p0?b4:b0))));
endmodule
