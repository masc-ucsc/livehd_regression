module expression_00153(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-5'sd11)!==(3'd5))>>((3'd6)==(5'sd12)))!==(5'd2 * ((3'd6)&(2'd2))));
  localparam [4:0] p1 = ({{(5'd9),(-5'sd9)},((-2'sd1)<=(5'd7))}>>{4{(4'd2)}});
  localparam [5:0] p2 = (4'd13);
  localparam signed [3:0] p3 = (({(-5'sd4),(2'd2),(4'd8)}<<{2{(4'd13)}})^~((3'd4)?(-5'sd10):(4'd7)));
  localparam signed [4:0] p4 = {1{{(!((4'sd4)^(5'd29))),{(5'd21),(4'sd6)}}}};
  localparam signed [5:0] p5 = (|({3{(3'd2)}}&&((3'sd1)^(4'sd4))));
  localparam [3:0] p6 = (4'd7);
  localparam [4:0] p7 = {1{{2{(~&(2'd0))}}}};
  localparam [5:0] p8 = ({2{(^(-2'sd0))}}>>(-(|((3'd7)===(3'sd2)))));
  localparam signed [3:0] p9 = ((|{3{(^(4'sd3))}})<<<(((2'd0)&&(-3'sd1))+((3'd0)+(2'sd1))));
  localparam signed [4:0] p10 = {((2'sd1)^~(5'sd14))};
  localparam signed [5:0] p11 = (({4{(2'sd1)}}&&(~&(-3'sd1)))?((&(5'sd10))?((-5'sd12)<<<(3'd2)):((4'd4)<(-5'sd10))):(((-4'sd2)?(4'd1):(4'd12))<(~^(3'sd2))));
  localparam [3:0] p12 = {2{(3'sd1)}};
  localparam [4:0] p13 = {1{{2{((5'd3)&&(-3'sd3))}}}};
  localparam [5:0] p14 = {1{(4'sd3)}};
  localparam signed [3:0] p15 = {(4'd10),(5'sd9)};
  localparam signed [4:0] p16 = {4{(4'sd7)}};
  localparam signed [5:0] p17 = (+(-5'sd2));

  assign y0 = (&(|((+(p0*p17))?((p11<p5)*(+p11)):(~(~(^p10))))));
  assign y1 = (+(((-(+p17))<=(p11>p6))|(!(-((a5^~a5)>=(-p3))))));
  assign y2 = (!{{((a1|b3))},((&b4)&&{p4}),{(b1?p3:b0)}});
  assign y3 = ((5'sd14)>>>$unsigned($signed(((p10^~b5)))));
  assign y4 = {2{(-3'sd0)}};
  assign y5 = ({4{(p15<p0)}}^(3'd2));
  assign y6 = (3'sd3);
  assign y7 = ((($unsigned(a1)<<<(b4!==b0))^$signed({b3,a1}))===(((6'd2 * b0)|{a1})!==((b5^~b0))));
  assign y8 = (((a2!==a4)^(~^b3))?((a5?p9:p16)^{p1,p7}):({a1}>>(4'd2 * p8)));
  assign y9 = (&(((^p10)?{p13,b1,p11}:(a3?a5:p4))?((~&p17)?(~|p6):(~|b5)):(~^{(p10?b3:a3),{a5,p13,p1}})));
  assign y10 = (((p8/p2)*(a0?p1:p16))<<((p16>>p12)^~(p7<<p6)));
  assign y11 = ({4{p0}}?(p9?p14:p15):(+p9));
  assign y12 = {p11,p6};
  assign y13 = ((((a3?a2:p13)?(b2+p0):(b5>=a5))-{(b3&&b3),(b1?p0:p15),(b5?a3:b3)})^(((p4<<p11)&&(a5|a5))||{1{((p7?p9:p6)=={2{b0}})}}));
  assign y14 = (2'sd1);
  assign y15 = (!((3'sd2)>>>(((p9%b1)<(b4?b3:a3))+((p16%p1)<(p10*a2)))));
  assign y16 = ({1{{2{(~^(p7?b0:b5))}}}}?{2{(!(p12?p0:p4))}}:{2{(p9==b5)}});
  assign y17 = (3'd3);
endmodule
