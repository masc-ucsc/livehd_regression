module expression_00150(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|((-4'sd2)?(5'd14):(5'd27)));
  localparam [4:0] p1 = (|{(^((2'd0)==(-4'sd5))),{2{(~&(5'sd4))}},{1{((2'd1)<<(5'sd15))}}});
  localparam [5:0] p2 = (((2'sd1)<=(4'd8))?((3'd4)?(5'd18):(-3'sd3)):((3'sd3)?(4'd5):(5'd9)));
  localparam signed [3:0] p3 = ((-(!(~&{1{(-3'sd0)}})))<(~(|((2'sd0)>>(-3'sd1)))));
  localparam signed [4:0] p4 = {2{(2'd3)}};
  localparam signed [5:0] p5 = (~(((2'sd0)?(2'd3):(5'd17))!={4{(5'd13)}}));
  localparam [3:0] p6 = {1{(~^(|((-3'sd2)>(-5'sd11))))}};
  localparam [4:0] p7 = {2{{2{(-2'sd0)}}}};
  localparam [5:0] p8 = {(2'd3),(2'sd1)};
  localparam signed [3:0] p9 = (((4'd11)+(2'd2))&&((5'd16)>>>(4'd4)));
  localparam signed [4:0] p10 = ((((-2'sd0)===(3'd1))?((-2'sd1)?(2'd0):(3'd0)):((2'sd0)?(2'd2):(3'd4)))<<<(4'd2 * ((4'd12)>(5'd6))));
  localparam signed [5:0] p11 = {{{((-2'sd1)<<(2'd0)),{2{(-3'sd0)}}}},{{(4'd7),(-2'sd1),(-5'sd4)},((3'sd1)?(4'd10):(5'sd13)),(2'sd0)}};
  localparam [3:0] p12 = ({{{(-5'sd7)}}}?((-3'sd0)?(2'sd0):(-3'sd3)):((4'sd3)?(5'sd4):(3'sd1)));
  localparam [4:0] p13 = ((((4'sd1)-(5'd20))^((5'sd5)<=(2'd1)))===({((5'd9)-(3'd7))}===((-5'sd9)^(3'd4))));
  localparam [5:0] p14 = (~((-4'sd1)&&(4'd5)));
  localparam signed [3:0] p15 = (~&(((2'd1)<<(4'd5))>((-2'sd0)?(2'd3):(2'd0))));
  localparam signed [4:0] p16 = (((2'd1)===(-2'sd0))?((-2'sd0)>>(4'd10)):((2'd2)^~(4'sd7)));
  localparam signed [5:0] p17 = {(((-3'sd3)===(4'd6))&&((3'd5)?(4'd14):(5'sd12))),{{(4'd14),(3'd5),(2'sd0)},{(2'd3),(5'd23),(3'sd0)}}};

  assign y0 = {3{(p15!=p4)}};
  assign y1 = (+((~^{((a0^~a5)=={1{a2}}),(~^{p1,a3,p13})})<={((-{3{a4}})!=={2{(a0&&a1)}})}));
  assign y2 = (^(((4'sd4)?(p15?p5:p8):(p1?p13:p8))<(-((&p13)?(p7*b1):(p16!=a3)))));
  assign y3 = (2'sd1);
  assign y4 = {{(~|(+(~&p9))),{$signed(p1),(~&p17)},{p7,p5,p17}}};
  assign y5 = $signed((|$unsigned(($signed((~|(^(~&p13))))))));
  assign y6 = (~|(^(2'sd0)));
  assign y7 = ((4'sd0)<={4{(p7+b2)}});
  assign y8 = (((p0!=p4)?(p8!=a5):(a3!=p9))?((4'd14)!==(b0?a2:a1)):(4'd2));
  assign y9 = ($unsigned($unsigned(p4))&{3{p15}});
  assign y10 = ((p9>>p13)!=(4'd2 * p6));
  assign y11 = (p13<=b4);
  assign y12 = {3{(-({2{{2{b4}}}}))}};
  assign y13 = ((b4?p13:p15)?{(a2?p11:p4)}:(b2?b2:a0));
  assign y14 = (2'd0);
  assign y15 = (-(~^(~^(~(4'sd5)))));
  assign y16 = (~&{2{(+(p7&p16))}});
  assign y17 = (~($unsigned((2'd0))*(p3+b0)));
endmodule
