module expression_00226(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((|(3'd2))^((-2'sd0)<<<(5'd16)));
  localparam [4:0] p1 = (((((3'd2)<<<(5'sd13))==((5'sd6)>(4'sd0)))<<{(5'd4),(2'd2),(2'd2)})!=((((4'd13)?(3'd2):(-2'sd0))>((5'd14)>>>(2'sd1)))-(3'd2)));
  localparam [5:0] p2 = (((~^(5'd22))?((2'd0)||(3'sd3)):((4'sd6)==(2'sd1)))<<(-(+((5'sd10)?(-2'sd1):(3'd1)))));
  localparam signed [3:0] p3 = (|{(3'd1),(-5'sd4),(3'd3)});
  localparam signed [4:0] p4 = (((-2'sd0)!==(3'd6))?(^(~(4'd7))):((2'd2)|(3'sd2)));
  localparam signed [5:0] p5 = ((5'sd6)|(3'sd2));
  localparam [3:0] p6 = {3{{2{(-3'sd1)}}}};
  localparam [4:0] p7 = {3{(&(2'd3))}};
  localparam [5:0] p8 = {2{(-3'sd0)}};
  localparam signed [3:0] p9 = (~((((-2'sd0)*(-2'sd0))>((5'd20)-(2'd3)))<<<(|(-(5'd2 * (2'd2))))));
  localparam signed [4:0] p10 = {(((4'd12)?(4'd8):(5'sd14))?((2'd0)<=(3'd3)):((5'd6)!==(-4'sd0))),(-2'sd0)};
  localparam signed [5:0] p11 = (6'd2 * (~|{3{(2'd0)}}));
  localparam [3:0] p12 = ({2{(2'd0)}}?{1{((-2'sd1)<<(5'd29))}}:((5'sd6)>>>(4'sd1)));
  localparam [4:0] p13 = ((3'd6)<<(-2'sd1));
  localparam [5:0] p14 = ((3'd4)-((4'd5)!==(5'd11)));
  localparam signed [3:0] p15 = ((((3'd3)^~(4'd1))>((-4'sd1)%(5'd30)))-(((-3'sd0)<(3'sd0))!==((2'sd1)|(-4'sd7))));
  localparam signed [4:0] p16 = (^(+{3{(^(~(-5'sd13)))}}));
  localparam signed [5:0] p17 = ((5'sd6)?{3{(3'd0)}}:((-4'sd4)!==(-4'sd2)));

  assign y0 = {4{({2{a2}}&&(b3&a3))}};
  assign y1 = ((b3)&&(b2^p2));
  assign y2 = $unsigned(($signed((p14/p2))%p9));
  assign y3 = ({3{(b3)}}===(^{3{{3{a4}}}}));
  assign y4 = {1{p6}};
  assign y5 = {(6'd2 * $unsigned((a5<<<p1)))};
  assign y6 = {({3{p7}}>=(3'sd2)),(((p0<=p8)<(a3!=a0))+{(4'd3),(2'd3)})};
  assign y7 = (~(|(((b1>>>a3))<=((^b5)))));
  assign y8 = (3'd1);
  assign y9 = (|(((~&p3)?{p2}:(~p6))?$unsigned((-{(4'd7)})):$unsigned((2'd1))));
  assign y10 = $unsigned(({2{{2{a4}}}}==={4{b4}}));
  assign y11 = {4{(~{1{(~|(|b2))}})}};
  assign y12 = (-(+(-3'sd2)));
  assign y13 = ((4'd14)?((p3*p0)>=(|b1)):((p4!=p1)>>(p16>p0)));
  assign y14 = ((-5'sd8)==={2{(4'd7)}});
  assign y15 = ((3'd5)^(4'd2 * {b1,b1,b0}));
  assign y16 = (({b2,b5,b1}?{a2,b4,p13}:(p15?a2:p1))?((~^b3)?{b2,p13,p8}:(p7?p4:a1)):(+(~^{(!(b2?b0:b5))})));
  assign y17 = (5'd29);
endmodule
