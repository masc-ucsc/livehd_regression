module expression_00198(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd2),(5'sd10),(3'd7)};
  localparam [4:0] p1 = (5'd15);
  localparam [5:0] p2 = (^({((2'sd1)+(2'd3)),(&(4'd3)),(!(-5'sd2))}!=(((3'd6)>>>(3'd1))^~(!((3'd4)<(2'd1))))));
  localparam signed [3:0] p3 = (!{(~|(-3'sd1)),{(2'sd1)}});
  localparam signed [4:0] p4 = {1{(2'sd1)}};
  localparam signed [5:0] p5 = ((&(-{((3'd5)?(5'sd1):(3'd2))}))?(5'sd10):(~&((-4'sd3)?(-3'sd1):(3'sd1))));
  localparam [3:0] p6 = (3'd0);
  localparam [4:0] p7 = ({3{(4'd13)}}?{(2'd1)}:{(4'd13),(-4'sd1),(5'd29)});
  localparam [5:0] p8 = {(4'sd0),(-2'sd0)};
  localparam signed [3:0] p9 = ((|(+(-(^((-5'sd5)?(3'd1):(-4'sd0))))))==={1{((2'd3)!==((4'd8)?(-2'sd0):(4'd0)))}});
  localparam signed [4:0] p10 = (-4'sd6);
  localparam signed [5:0] p11 = ((4'd10)>>(~((5'sd11)<=(-3'sd0))));
  localparam [3:0] p12 = ((((3'sd1)<<(5'd7))&&((3'd4)?(4'sd5):(-2'sd1)))>>{3{((2'd3)===(5'd3))}});
  localparam [4:0] p13 = (|((((3'd4)&&(5'd24))>>>((3'd4)-(3'd5)))+{2{(&(2'd0))}}));
  localparam [5:0] p14 = {{(~^((3'd1)>=(4'd13))),(~|((-5'sd9)>>>(3'sd0)))}};
  localparam signed [3:0] p15 = (+(|((-2'sd1)<=(3'sd0))));
  localparam signed [4:0] p16 = ((((-4'sd1)?(2'd2):(2'd2))&&((4'd0)&&(-5'sd9)))>>>(((-5'sd14)&(-4'sd7))?((3'd5)!==(5'd25)):((3'd2)<<<(2'sd0))));
  localparam signed [5:0] p17 = {{(~|((&(~^(-4'sd3)))!=(~|((5'd3)+(4'd6))))),({2{(4'sd0)}}-(5'd2 * (3'd2)))}};

  assign y0 = (+{4{p13}});
  assign y1 = ((-3'sd2)?(a2^p16):(a0?p2:b2));
  assign y2 = (&($unsigned($signed((|((a0?b4:a0)^~(a1<b1)))))==={$signed({$unsigned((a4?a5:a3)),(a4?a5:b4)})}));
  assign y3 = ($signed(b0)?(~^a0):(-a1));
  assign y4 = (+(+(b1?a3:b3)));
  assign y5 = {1{({(3'd7),(p2<=a4),(~&p8)}<={2{(~&(p14&b3))}})}};
  assign y6 = ({({p15}?$unsigned(a1):(p7?p9:p0)),$signed((2'd1))});
  assign y7 = {{1{({3{b0}}^{p15,a3,a0})}},((a3&b0)!==(a5&a4))};
  assign y8 = (+(!(~&(~|{(5'd28)}))));
  assign y9 = ((5'd2 * (p14!=p12))<<<(((p2-p11)?(p13>>>p12):(~|p6))>>>(&((p12?p5:p1)<<(p11*p4)))));
  assign y10 = {{{a4,p16,b5},$unsigned((3'sd3)),(3'd5)}};
  assign y11 = $signed((+((a5===b1)*$unsigned((~^p12)))));
  assign y12 = (5'd31);
  assign y13 = ((((b5>>>a4)<(5'd2 * b0))===((a3<=b3)>(b5<a4)))===(((a4|a4)>=(b4!=b3))<<<((b5^~b1)<(b0===a1))));
  assign y14 = $unsigned(($signed($signed((p14/p12)))>=(&((p1!=p1)<=(p15?a0:p11)))));
  assign y15 = ((p3?b5:p13)?(p16?p12:p15):(p11|p1));
  assign y16 = $unsigned($signed(({4{($signed(a5)===(a0&b1))}})));
  assign y17 = (~&(b5|p5));
endmodule
