module expression_00932(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd1);
  localparam [4:0] p1 = ((3'sd2)<<(5'd2));
  localparam [5:0] p2 = ((+((2'd0)<(3'd7)))>((2'd1)>(-4'sd4)));
  localparam signed [3:0] p3 = (~^((((-5'sd7)^~(-4'sd6))^~(&(3'd3)))<<<(6'd2 * (3'd4))));
  localparam signed [4:0] p4 = (((-2'sd0)?(-3'sd3):(3'd5))?((2'd3)?(2'd1):(5'd16)):((-5'sd6)?(5'sd8):(4'sd0)));
  localparam signed [5:0] p5 = (-2'sd1);
  localparam [3:0] p6 = (((5'd31)>>(3'sd3))-((3'd3)^~(5'sd11)));
  localparam [4:0] p7 = ((({(4'd7),(-3'sd3)}^{(3'sd1),(5'd12),(-2'sd0)})<((3'sd2)?(5'sd0):(3'd6)))&&({1{(~&(~^(4'd8)))}}!==(!{(~|(-2'sd1))})));
  localparam [5:0] p8 = ({(+((4'sd6)>(2'd0))),((4'sd2)==(3'sd0))}^~(|{(~^((2'd1)!=(4'd0)))}));
  localparam signed [3:0] p9 = (&(|(-4'sd6)));
  localparam signed [4:0] p10 = ({((-2'sd0)>>(2'd0)),{4{(3'sd0)}}}>>({(-3'sd1),(2'd3)}<(-4'sd7)));
  localparam signed [5:0] p11 = {4{((-5'sd9)!=(4'sd0))}};
  localparam [3:0] p12 = {((!(!(4'd11)))||((4'd7)?(3'd3):(2'd3))),{({(3'sd2),(3'd3)}===(+((2'sd0)!==(-5'sd4))))}};
  localparam [4:0] p13 = {2{(5'sd14)}};
  localparam [5:0] p14 = (~|(-(4'sd2)));
  localparam signed [3:0] p15 = {4{(^(5'd5))}};
  localparam signed [4:0] p16 = {2{{4{(2'd3)}}}};
  localparam signed [5:0] p17 = {(((3'd5)+(3'd2))||((4'd9)^~(5'sd8))),((5'd7)&&(6'd2 * (5'd28)))};

  assign y0 = {4{(~&p6)}};
  assign y1 = ((((4'd14)^~(b1<=p16))<<(3'd1))|(3'd3));
  assign y2 = (5'd9);
  assign y3 = ((5'd2 * {2{p12}}));
  assign y4 = {4{(~|$signed({4{p11}}))}};
  assign y5 = {2{{3{(a4&&p16)}}}};
  assign y6 = (((((a5?a1:b5)==(a3?b1:b3)))+((a4?a3:b2)?(a0&&a2):$signed(a2)))!==((a5?b2:b5)*(a4?a3:b4)));
  assign y7 = (^b2);
  assign y8 = ((({2{a0}}>=(3'sd1)))<(5'd16));
  assign y9 = {(-5'sd6)};
  assign y10 = {1{{({1{p9}}?(b2&&p3):{4{p6}}),((p10^~a3)<{p7,a4})}}};
  assign y11 = {{{b1},(a3^a1),(b1&a2)},((a4|b0)&(p16>>>b2)),((b4?a2:a1)+(a0?b0:a2))};
  assign y12 = ((((2'd2)/b4)+($unsigned((a2||a1))%b4)));
  assign y13 = ((~^((p3^a2)?(p2?a0:p3):{p14,p3}))<<(-{(p1<=p11),(p2?p5:b5),{p8,p3,b2}}));
  assign y14 = (-$unsigned(p8));
  assign y15 = ((p0?p0:p11));
  assign y16 = {(+(a1>>>p16)),(-(~&p14)),{a0,a4}};
  assign y17 = {((b5<<<b0)>>>(5'd2 * a2)),(~&((p10>>>a5)-(b0<p9)))};
endmodule
