module expression_00611(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd20);
  localparam [4:0] p1 = (~&(|(4'd3)));
  localparam [5:0] p2 = (~|(~|(~&{3{(-4'sd5)}})));
  localparam signed [3:0] p3 = ((((4'd6)>>>(4'd10))==((-4'sd6)>(3'd1)))^(((-4'sd1)&(-5'sd8))<((-2'sd0)&(-2'sd1))));
  localparam signed [4:0] p4 = {4{(~((4'sd6)<=(3'd0)))}};
  localparam signed [5:0] p5 = (~^(~(-{2{((4'd5)?(5'd3):(2'sd0))}})));
  localparam [3:0] p6 = (((~&((-2'sd1)&(-3'sd2)))!=((2'sd1)>=(2'd2)))+(&(((-3'sd3)>(2'd2))>((3'd5)>>(5'd10)))));
  localparam [4:0] p7 = (({(4'd5),(5'd27),(2'd2)}&&((5'd1)^~(3'sd2)))<<<((~|((-5'sd2)==(-3'sd2)))!==((4'sd2)===(-4'sd7))));
  localparam [5:0] p8 = ((((5'sd1)||(-4'sd3))^~(~&(2'd2)))?(!(-(~|((2'd3)==(5'sd13))))):((~(3'sd2))+((3'sd2)>(4'd11))));
  localparam signed [3:0] p9 = (~|((~|(3'd0))==={2{(-5'sd8)}}));
  localparam signed [4:0] p10 = (3'sd2);
  localparam signed [5:0] p11 = (-{((5'sd13)|(4'sd3))});
  localparam [3:0] p12 = ({(4'sd5),(4'd4)}?(+(-3'sd0)):((-3'sd3)?(3'd2):(-2'sd1)));
  localparam [4:0] p13 = {1{{4{(3'd4)}}}};
  localparam [5:0] p14 = {(-5'sd13),(4'sd5)};
  localparam signed [3:0] p15 = (|(-5'sd13));
  localparam signed [4:0] p16 = (+((5'd2 * (5'd28))?(-2'sd1):((-5'sd8)?(-2'sd1):(-5'sd10))));
  localparam signed [5:0] p17 = (-4'sd7);

  assign y0 = {(b3?b2:p13),(|(a5?p5:p11))};
  assign y1 = ({4{(b5===a1)}}<((p12?p14:b3)^(5'd2 * p0)));
  assign y2 = (-((p6<=p0)&&(a1===b2)));
  assign y3 = {3{(~b4)}};
  assign y4 = {2{{1{{4{b4}}}}}};
  assign y5 = (~|(|(-3'sd1)));
  assign y6 = {{(^(-(&p0))),({a4,p17})},{{{b2,b4},{b4}},{(^b5),$unsigned(a4)}}};
  assign y7 = (((~^p10)?(p3&&a2):{2{p2}})?(2'sd1):{1{{2{$unsigned(p14)}}}});
  assign y8 = (((!p5)^~(p17^~p7))?((b1?p13:p5)<=(b0?p8:a3)):(~&((-2'sd1))));
  assign y9 = (((p16?p7:p9)?(p3?a0:p14):(p13?p5:b0))?((a4?p2:p3)?(a1?p7:p16):(p3?p6:p11)):((p4?p15:p12)?(p11?p8:p15):(b5?a3:p7)));
  assign y10 = (4'sd3);
  assign y11 = ((!(~^(3'sd3)))?(5'd17):(~^{2{p16}}));
  assign y12 = (b4!==b0);
  assign y13 = (((p10?p17:p9)&(p16>=p3))?((b4&p1)>>(p16==p3)):(a2?p0:p10));
  assign y14 = (&(3'd3));
  assign y15 = (!a3);
  assign y16 = {1{{3{(|{4{p15}})}}}};
  assign y17 = $signed({(({a0})?(a0<b0):$signed((3'd3))),((2'd2)^(b4?b4:b2))});
endmodule
