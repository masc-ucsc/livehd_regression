module expression_00132(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd0)===(-3'sd2));
  localparam [4:0] p1 = (5'd8);
  localparam [5:0] p2 = (~|(^(((3'd6)?(-3'sd0):(5'd3))?((2'd2)?(3'sd0):(3'd4)):(5'd2 * (2'd0)))));
  localparam signed [3:0] p3 = (-((((3'd0)>>(5'd25))|(^(-5'sd6)))==(((-2'sd1)<(3'd6))||(~^(3'sd0)))));
  localparam signed [4:0] p4 = ((({1{(3'd5)}}<={3{(2'd1)}})<<<{3{(3'd2)}})>>>(3'sd0));
  localparam signed [5:0] p5 = (~|(4'sd1));
  localparam [3:0] p6 = ((((5'sd13)?(5'd17):(-3'sd3))?((-4'sd7)<<(-4'sd1)):((5'd12)!=(2'd3)))<({2{(2'sd1)}}<=(3'd5)));
  localparam [4:0] p7 = (((-3'sd2)?(-4'sd4):(-5'sd9))?{(-4'sd6),(2'sd0),(2'd2)}:((-5'sd14)?(2'sd0):(-2'sd0)));
  localparam [5:0] p8 = (4'sd5);
  localparam signed [3:0] p9 = (-(&{4{{1{{3{(4'sd6)}}}}}}));
  localparam signed [4:0] p10 = {4{(-(-2'sd0))}};
  localparam signed [5:0] p11 = {3{{(5'd10),{3{(3'd4)}}}}};
  localparam [3:0] p12 = (5'd20);
  localparam [4:0] p13 = {{{{(3'd0),(2'd1),(2'd0)},(-(2'd0))},{{(-5'sd4)},{(3'sd2)}}},{(2'd3)}};
  localparam [5:0] p14 = {{2{(3'd5)}}};
  localparam signed [3:0] p15 = (!(((!(3'd1))?(-(5'sd8)):((5'sd6)?(2'd1):(-5'sd5)))<(~|(((-2'sd1)&&(-2'sd0))?((4'd8)>(-3'sd0)):((5'd30)>>>(-4'sd2))))));
  localparam signed [4:0] p16 = (((~&(2'sd0))^{4{(4'd9)}})||(((4'd8)>(3'd3))===((5'd2)<(-5'sd5))));
  localparam signed [5:0] p17 = (~|((!(5'sd3))!=((-4'sd2)||(-4'sd6))));

  assign y0 = {$signed($signed(p7)),(b0===a0),((p10<<a2))};
  assign y1 = (-3'sd3);
  assign y2 = ({(-{b3})}>>(!(~&(p1<<b5))));
  assign y3 = {2{{(2'sd0)}}};
  assign y4 = ({3{(p11>=p6)}}>{{2{{1{a4}}}},(-(p2?p6:p9))});
  assign y5 = ((5'sd3)?(-2'sd1):(p10?b5:a0));
  assign y6 = (!$unsigned((((3'd7)>=$unsigned((p13!=p6))))));
  assign y7 = (-b5);
  assign y8 = (({4{b2}}>>{3{b4}})?(&((~p15)>=(b2>=p17))):((p1||a4)<{4{a2}}));
  assign y9 = (~&(((6'd2 * a0)>>(a4+p12))<=((p8<<p11)<<(b0%b5))));
  assign y10 = ((+(4'd8))?((a1>a2)==={b4,a4}):((2'd3)^~(5'd28)));
  assign y11 = (a5);
  assign y12 = ((((b1^a3)<{1{b1}})!=={4{a1}})!=(((a1!==b5)-(p17&b5))^~{(b1<<<p10)}));
  assign y13 = {($signed(p0)?(^b0):(b5?p1:a3)),((b0?a0:b3)|$signed(a3))};
  assign y14 = (a5>=p14);
  assign y15 = (&(({a5,a4,a0}?{3{b5}}:(b3?b2:a5))^~(~|((~&(a0?a0:b4))?(a2>p0):(!(b0?p9:b3))))));
  assign y16 = (+(2'd1));
  assign y17 = (((b0>a0)>(a4!=b0))?((p4>b0)>=(p7|b4)):((a1<=b3)!==(b2==a4)));
endmodule
