module expression_00208(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^((+(+{((4'sd2)!==(4'd4)),{(-4'sd2),(4'd15),(2'd1)},((3'd2)<<(3'd4))}))>>(6'd2 * ((3'd1)^~(2'd1)))));
  localparam [4:0] p1 = (3'd0);
  localparam [5:0] p2 = {2{(~|((~|((-2'sd1)&(4'sd4)))^((2'sd0)-(4'sd3))))}};
  localparam signed [3:0] p3 = (({(2'sd1),(5'sd14),(-3'sd2)}&(6'd2 * (3'd2)))!==(~{(+{(+(~&(-5'sd7)))})}));
  localparam signed [4:0] p4 = (4'd3);
  localparam signed [5:0] p5 = (-(^(&{((2'sd1)<(5'd24)),((5'd28)<<<(-5'sd4))})));
  localparam [3:0] p6 = (~((4'd11)?(2'd3):(2'sd0)));
  localparam [4:0] p7 = ((&(5'sd13))<(|(5'd26)));
  localparam [5:0] p8 = (((5'd4)>(-3'sd3))!=((-2'sd1)?(2'd0):(-3'sd1)));
  localparam signed [3:0] p9 = (~(2'sd1));
  localparam signed [4:0] p10 = ((((3'sd2)+(3'd6))|((4'sd2)&(3'd4)))&{3{((-5'sd1)<=(3'd5))}});
  localparam signed [5:0] p11 = ((-2'sd1)?(5'd16):(-5'sd1));
  localparam [3:0] p12 = (-((^((3'd4)?(-3'sd1):(5'd24)))?(~^(~^((5'd31)?(3'd0):(4'sd6)))):((5'd3)?(4'd3):(4'd6))));
  localparam [4:0] p13 = (~{(+{(~^{(+(+(-2'sd0)))}),(~{{{(5'd21),(3'sd1),(4'd9)}}})})});
  localparam [5:0] p14 = (~|(!{(~(~(4'd15))),(&{(3'sd2),(2'd0)}),{(-2'sd1),(2'd3)}}));
  localparam signed [3:0] p15 = (((2'd3)|(-4'sd5))*(2'sd0));
  localparam signed [4:0] p16 = (((2'd3)<=(5'sd14))||((-5'sd12)+(4'd13)));
  localparam signed [5:0] p17 = ((4'd3)+(-5'sd14));

  assign y0 = (~&(a0));
  assign y1 = {2{p2}};
  assign y2 = (!(|(~&p15)));
  assign y3 = (4'd2 * (3'd2));
  assign y4 = (3'sd3);
  assign y5 = ((&(&$unsigned(((!(~&(~^(~^$signed(p17)))))||((~(p15<<p10))!=(|(p11>>p9))))))));
  assign y6 = (5'sd10);
  assign y7 = (5'd16);
  assign y8 = (a4>>b3);
  assign y9 = (((~|(-((4'd2 * b0)<=(a0==p16)))))-(((p6)||(a5>>a3))^~{p13,b1,p13}));
  assign y10 = (a0>=p16);
  assign y11 = (p3-b1);
  assign y12 = ((({a0,b1}===(a4&&a3))+(p13?p16:p10))^(((p12+p0)|(p9||p16))!=((p12?p2:p3)<=(p0<<p0))));
  assign y13 = ({(~^p10),(b5?p2:b3),(~&p9)}!=((b2?p1:a3)?(p11?p2:p7):(a4!==a5)));
  assign y14 = (($unsigned(((a4<=b1)<<(5'd14))))-{1{(3'd1)}});
  assign y15 = (!(&(3'd2)));
  assign y16 = (5'sd10);
  assign y17 = {3{$signed((!{2{{2{p0}}}}))}};
endmodule
