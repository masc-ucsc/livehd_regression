module expression_00957(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{{3{((3'd2)?(5'd17):(-4'sd6))}}}};
  localparam [4:0] p1 = (!(((~(3'd1))===((3'd1)&(2'sd1)))||((&(2'd1))>>>{(4'd8),(3'sd3)})));
  localparam [5:0] p2 = ((((3'd3)?(2'sd1):(5'd5))?((4'd12)>>(2'd2)):{3{(2'sd0)}})<(|({(5'sd8),(4'd6),(2'd0)}||{3{(3'd0)}})));
  localparam signed [3:0] p3 = ((((5'd17)+(2'd1))<<<(3'd4))&&(-3'sd1));
  localparam signed [4:0] p4 = {(3'sd2)};
  localparam signed [5:0] p5 = {((4'sd4)-(-3'sd0)),(-(5'sd12))};
  localparam [3:0] p6 = (!(-3'sd1));
  localparam [4:0] p7 = (~|((~&(+(~&(-(&((3'd7)<(2'd3)))))))<<<(|(|(~^((+(3'd4))<(|(4'sd0))))))));
  localparam [5:0] p8 = (~(-2'sd0));
  localparam signed [3:0] p9 = (({1{{4{(4'sd6)}}}}?((-2'sd1)>>(4'd5)):((4'd5)?(2'd1):(2'sd1)))||{2{((4'd6)?(4'd1):(4'd9))}});
  localparam signed [4:0] p10 = (2'd2);
  localparam signed [5:0] p11 = (2'd1);
  localparam [3:0] p12 = (((4'd10)<=(-3'sd3))|((2'd2)||(4'sd6)));
  localparam [4:0] p13 = ((~^{2{(2'd3)}})!==((2'd2)^(-5'sd14)));
  localparam [5:0] p14 = (+(5'd4));
  localparam signed [3:0] p15 = (~^{{(3'd3),{(5'd27)},(~|(3'sd3))}});
  localparam signed [4:0] p16 = (((4'sd5)?(2'd2):(-4'sd7))>=((3'sd1)===(4'd0)));
  localparam signed [5:0] p17 = ((&(((-5'sd6)-(2'd1))>((3'sd3)?(3'd0):(-5'sd10))))^(((4'sd4)|(-3'sd2))<<<(5'd30)));

  assign y0 = {4{{1{p7}}}};
  assign y1 = ((p16&&a2)<<<(p13&&p6));
  assign y2 = ($unsigned(((~b3)===(6'd2 * b0)))?((b1|b0)===(a3<<a1)):(5'd2 * (b0?a0:p12)));
  assign y3 = {{(3'd5),{((a4|a1)==(|(a3<p7)))},(3'sd2)}};
  assign y4 = ((p7)>>(b5!==a3));
  assign y5 = (2'sd1);
  assign y6 = ((~^((2'sd1)==$signed((5'sd13)))));
  assign y7 = ((p17^b3)^~(a4===a1));
  assign y8 = ({4{(+a3)}}<=((p0?p11:p9)?(a5?p10:p5):(p12<=p10)));
  assign y9 = (+(-(~(2'd2))));
  assign y10 = ((b3?a4:p6)?(a5?b5:a0):{4{b5}});
  assign y11 = {1{{{(p13<=a0),(a2|p12)}}}};
  assign y12 = {{($signed({a3})),(~^(a0^~b2))},((~|(a4))?$signed($signed(a5)):(b0?a5:p7))};
  assign y13 = ((3'd6)?((p2>p4)&&{1{a0}}):(3'd2));
  assign y14 = (!(3'd1));
  assign y15 = {4{(~&{1{p1}})}};
  assign y16 = (~&(~&(&(-p6))));
  assign y17 = {(2'd1),((p0?p6:p0)>(p9<p6)),{(2'd1),(p9?p14:p3)}};
endmodule
