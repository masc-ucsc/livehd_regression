module expression_00140(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((5'd8)&&(3'd7))&&((5'd20)===(4'd6)))^(((4'd14)<<<(-3'sd1))>>((-2'sd0)===(3'd4))));
  localparam [4:0] p1 = ((5'd17)>=(-3'sd3));
  localparam [5:0] p2 = ((3'd7)?(5'sd1):(-2'sd0));
  localparam signed [3:0] p3 = ((3'd4)?(2'd0):(5'd29));
  localparam signed [4:0] p4 = (&{1{((~&(2'sd0))+(+(4'd2)))}});
  localparam signed [5:0] p5 = ((-4'sd4)?(4'd2):(5'sd15));
  localparam [3:0] p6 = (((3'd1)^(4'd9))?((3'd6)|(5'd2)):(~^{2{(4'd0)}}));
  localparam [4:0] p7 = (~|{4{{4{(5'd15)}}}});
  localparam [5:0] p8 = (|(~|(^(~^(~^(4'd2 * ((4'd10)>(2'd1))))))));
  localparam signed [3:0] p9 = ({(-2'sd0),(5'd7),(-5'sd6)}?{(4'd3),(3'd7),(5'd13)}:((2'sd0)==(-3'sd2)));
  localparam signed [4:0] p10 = (((-5'sd9)^(5'd0))>=((2'd0)>(4'd0)));
  localparam signed [5:0] p11 = (-3'sd0);
  localparam [3:0] p12 = {1{((+(2'd0))&&{2{(4'sd4)}})}};
  localparam [4:0] p13 = (2'sd0);
  localparam [5:0] p14 = ((((3'd3)?(5'sd15):(3'sd1))<<((2'sd1)?(5'd7):(2'sd1)))>>>(4'd0));
  localparam signed [3:0] p15 = (-((3'd4)<<(-5'sd15)));
  localparam signed [4:0] p16 = {(-4'sd0),(3'd4)};
  localparam signed [5:0] p17 = ((3'd6)&&(-4'sd3));

  assign y0 = {2{{2{{1{{1{b3}}}}}}}};
  assign y1 = {3{(+{{a4,b0,b1}})}};
  assign y2 = {{3{a4}}};
  assign y3 = (((((b0)<<(b3^p15)))|$signed(((b3>=a2)^~(|p9))))!=($unsigned((~((~|b1))))<((~|a0)<=(b3<=a1))));
  assign y4 = $unsigned((2'd3));
  assign y5 = (^((|{$unsigned((~&({p15}))),(|(!{(|p6)})),(-(~{{2{p11}}}))})));
  assign y6 = {2{{(p14?a1:b4),(~|p14),(p1?p11:p8)}}};
  assign y7 = {{$signed((($signed(b1)<$signed(a1))===({a2,b2}>>$signed(b4))))},($unsigned(({$signed(b4)}))&{(b3),$signed(b3),(p7|p7)})};
  assign y8 = (3'd2);
  assign y9 = {2{(^(^{(b4>b0)}))}};
  assign y10 = (a2-a0);
  assign y11 = (~^(a0-p10));
  assign y12 = {({4{p3}}?{a0}:{4{a0}}),(3'd0)};
  assign y13 = (!((((p15/p9)?(p5?p9:p1):(p8%p12))>>>((p3>=p14)|(p15<p12)))));
  assign y14 = {3{{2{((p2))}}}};
  assign y15 = ((({b0,a1,b3}&&{b1,a4})!=(|{{4{b2}}}))||({(b2<<a3)}!=({p6,p8}>>(-p4))));
  assign y16 = ((2'd0)!=$signed((~|(^p10))));
  assign y17 = (~^(~&(({p0,p14,a2}?{4{p15}}:{p17})?{{p5},(p2?p16:p14),(p8?p1:p1)}:{(^{p7,p3})})));
endmodule
