module expression_00898(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(-((+((-(-3'sd2))<<<((-2'sd0)>=(-5'sd1))))|(((-5'sd12)|(3'd3))?(~(3'sd1)):((5'd24)?(5'd19):(3'd3))))));
  localparam [4:0] p1 = ((((5'd4)?(2'sd1):(-2'sd1))?((2'd1)?(4'sd1):(4'd15)):((-4'sd6)?(4'd9):(3'sd2)))?{2{(|(5'd5))}}:(((5'd28)^~(-2'sd0))>>{4{(5'sd14)}}));
  localparam [5:0] p2 = ((((2'sd1)+(-3'sd3))?(+(3'd5)):{3{(2'd2)}})&&((~^(-5'sd4))&&{4{(-5'sd13)}}));
  localparam signed [3:0] p3 = ({((5'd31)-(-2'sd1)),{4{(2'sd1)}},{(2'd1)}}^{{3{(3'd5)}},{(3'd0),(-4'sd0),(5'd26)}});
  localparam signed [4:0] p4 = ((^(!(-(3'd1))))>={((~^(~&(4'sd6)))!=((5'sd7)&&(3'd0)))});
  localparam signed [5:0] p5 = (3'sd1);
  localparam [3:0] p6 = ((5'd20)&&(-3'sd2));
  localparam [4:0] p7 = (((4'd15)?(2'sd1):(4'sd0))?((4'sd2)?(-3'sd0):(5'd18)):(((4'sd1)?(2'd2):(-4'sd0))&((-3'sd0)?(-2'sd0):(3'sd3))));
  localparam [5:0] p8 = (((4'd2)-(-2'sd1))==(|((-4'sd0)<<(-5'sd12))));
  localparam signed [3:0] p9 = ((&((-3'sd1)>=(2'd0)))>>((-5'sd4)==(5'sd6)));
  localparam signed [4:0] p10 = ((-2'sd1)|(2'sd1));
  localparam signed [5:0] p11 = (!(-5'sd3));
  localparam [3:0] p12 = (|(((|(^(5'sd5)))^((2'sd1)!=(5'd21)))|(5'd2 * (+{(3'd6),(3'd1)}))));
  localparam [4:0] p13 = ((^((5'sd14)<(3'd3)))?(~&(-2'sd0)):(~^(3'd4)));
  localparam [5:0] p14 = {{{3{{(-3'sd2),(-5'sd10),(5'sd2)}}}},(4'sd4)};
  localparam signed [3:0] p15 = ((((5'd7)?(5'd10):(-3'sd0))?{(2'sd0)}:{(5'sd8),(3'd6)})?{((-5'sd15)?(5'd2):(4'd14))}:(-2'sd0));
  localparam signed [4:0] p16 = (((3'd3)|(5'sd9))>>((4'd4)*(4'd8)));
  localparam signed [5:0] p17 = (^(~(~&{{4{(3'd4)}},(((2'sd0)^(5'd12))!=(~^(-2'sd0)))})));

  assign y0 = {({{1{{$signed($signed(a4)),{2{p6}},{a3,p9}}}},$signed({{4{p7}},(-{p1,p6}),$signed({1{p16}})})})};
  assign y1 = (&({{p1,p5,p2}}?(&(p3|b3)):(p5?p7:p1)));
  assign y2 = (p3?p10:p13);
  assign y3 = (~|((~(5'sd8))));
  assign y4 = (~&(3'd7));
  assign y5 = {{((!p4)+{p8,p14}),((~^p12)>>>{p14}),((|p15)&&(&p8))}};
  assign y6 = (~&(!a3));
  assign y7 = {3{p6}};
  assign y8 = ((&((~(a4!==b4))|(-(p2<=p7))))>({(b3<<<p15)}&&(p2<<<b0)));
  assign y9 = ({{2{{a2}}},({b3,p11,b5}),{1{{{3{p15}},(b5)}}}});
  assign y10 = ((p0>>p0)^$signed((a3%p2)));
  assign y11 = ((~p9)||(b3&&p7));
  assign y12 = (|a5);
  assign y13 = $signed((|(-(($unsigned((b4+a4))===$unsigned((+a5)))<<<((a1<<p5)?$signed(b3):$unsigned(p6))))));
  assign y14 = ((^{a3})?(^(2'd0)):(a1===a0));
  assign y15 = ({3{{{(a3)},(~^(&a3))}}});
  assign y16 = (5'd11);
  assign y17 = (~&(b0^~b2));
endmodule
