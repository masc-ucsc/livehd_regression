module expression_00565(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(^(~|(~&(4'd2)))));
  localparam [4:0] p1 = {2{(3'sd2)}};
  localparam [5:0] p2 = {{(6'd2 * ((3'd7)?(4'd3):(2'd0)))},(((4'sd1)?(4'sd0):(5'd15))||((-2'sd0)?(-5'sd15):(5'd2)))};
  localparam signed [3:0] p3 = ((4'd12)||(3'd4));
  localparam signed [4:0] p4 = (~&(3'd3));
  localparam signed [5:0] p5 = ({4{{2{(-3'sd2)}}}}>>(|(~&{1{(((5'd13)&(3'd7))^(4'sd6))}})));
  localparam [3:0] p6 = {(((3'd2)<<<(-3'sd1))>>>((-4'sd4)===(4'sd1))),(((2'd0)||(3'd0))!=={(5'd3)}),{({(3'd2),(3'd5),(2'd0)}>>{(-4'sd5),(-2'sd1),(2'sd0)})}};
  localparam [4:0] p7 = (^(~({2{((3'd3)===(3'd3))}}?(((5'd10)<(5'd8))<<<(+(-4'sd3))):{1{((5'sd2)>(4'd6))}})));
  localparam [5:0] p8 = {1{({{1{{(4'd8),(3'sd0)}}},(4'd2 * (5'd26))}<<<{2{{(3'sd2),(3'd1),(4'sd1)}}})}};
  localparam signed [3:0] p9 = ((((5'd21)-(3'sd3))!=((-4'sd7)^~(-4'sd6)))!==(4'd2 * ((3'd0)!=(2'd2))));
  localparam signed [4:0] p10 = ((((2'd1)^~(-2'sd0))<=((-2'sd0)*(2'd0)))===(((5'd31)?(2'sd0):(2'd3))==((3'sd3)<=(-5'sd6))));
  localparam signed [5:0] p11 = {4{{{4{(5'sd10)}}}}};
  localparam [3:0] p12 = ((((2'sd0)?(-5'sd7):(3'd6))%(4'd12))>>>(((-2'sd0)?(-2'sd1):(-4'sd3))!=(+(-5'sd11))));
  localparam [4:0] p13 = (-(~|(|{3{(5'd1)}})));
  localparam [5:0] p14 = (&(4'd2));
  localparam signed [3:0] p15 = ((^(&(3'd5)))<((5'd16)^~(4'd13)));
  localparam signed [4:0] p16 = (((+((3'd1)?(3'sd1):(3'd2)))?((2'd3)+(-2'sd1)):((4'd15)+(4'd13)))>>(((-2'sd1)^(3'd3))?{(2'd2),(4'd15),(5'd12)}:((-3'sd0)==(5'd9))));
  localparam signed [5:0] p17 = {1{{1{({2{{(~^(4'sd5))}}}<<{2{{1{(-(2'd3))}}}})}}}};

  assign y0 = ((~^(~p10))>>{p10,p14,b3});
  assign y1 = (~|(|(^a2)));
  assign y2 = (&{b4,p2,a3});
  assign y3 = {1{{4{{{b5,p0,a0},{2{b5}},{3{a3}}}}}}};
  assign y4 = (+(((~p3)^~(p3*a4))?(-5'sd1):$unsigned((5'sd6))));
  assign y5 = ({1{(|((&b5)?(~&p2):(2'sd1)))}}|{1{{1{({4{a3}}?(a4>>b0):(b3?a3:p6))}}}});
  assign y6 = {{{p4},(b0|p10)},((a2>=b4)&(p17+a4))};
  assign y7 = ((~&(-p1))+(b2>>b0));
  assign y8 = (~(3'd5));
  assign y9 = ((((a2===b3)*(b5&&a4))||((a4*a4)<=(p11&p14)))!=(((-b2)*(p13<p17))^~((a1|a1)<<(a0==p11))));
  assign y10 = (~|(&p14));
  assign y11 = (({$signed({p6,a0,b0})})<(({p3,a1})<=$signed((4'sd7))));
  assign y12 = (~^{1{a3}});
  assign y13 = (p14>=a3);
  assign y14 = {3{(a2?a4:b2)}};
  assign y15 = ({p8,p7,a3}+{2{p14}});
  assign y16 = {b4};
  assign y17 = ($signed((((~(p4>p17)))==(~|(a4!=a5))))>=$signed((^((&(!a1))-(!(~&b4))))));
endmodule
