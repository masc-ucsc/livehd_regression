module expression_00423(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd0);
  localparam [4:0] p1 = {2{(~^(2'd2))}};
  localparam [5:0] p2 = (((&(4'sd7))||((2'sd1)<(2'd1)))&{3{(5'd21)}});
  localparam signed [3:0] p3 = ((((-3'sd1)&&(4'd15))==((-2'sd0)<<(2'sd0)))&(((5'sd3)<<<(4'sd0))?((4'd3)||(-5'sd4)):((3'sd1)|(4'sd0))));
  localparam signed [4:0] p4 = {{((2'sd1)>=(3'd7)),((2'sd1)-(4'sd2)),{(4'd8)}}};
  localparam signed [5:0] p5 = ((5'sd2)?(-2'sd0):(-5'sd6));
  localparam [3:0] p6 = (6'd2 * ((2'd0)^(4'd2)));
  localparam [4:0] p7 = ((4'd9)>(3'd6));
  localparam [5:0] p8 = {((-2'sd0)?(5'd8):(-2'sd1)),((4'd10)?(-5'sd3):(3'sd2)),({(3'd2)}||((4'sd2)?(4'd6):(2'd3)))};
  localparam signed [3:0] p9 = ({{(5'sd6),(3'd5),(4'd13)},((2'sd0)+(4'd4))}||{{((5'd12)>>(5'd2))}});
  localparam signed [4:0] p10 = (((~|((4'd10)-(-4'sd3)))<<((2'sd1)==(3'd0)))>>{((5'd31)-(5'd15)),((2'd2)?(5'sd6):(5'd27)),(+(-5'sd10))});
  localparam signed [5:0] p11 = (-2'sd0);
  localparam [3:0] p12 = (4'd6);
  localparam [4:0] p13 = (~&(~&((4'sd0)?(4'sd0):(5'd29))));
  localparam [5:0] p14 = (~^(~&(+(~&((~^((-3'sd1)%(5'd9)))<=(^(+(-5'sd4))))))));
  localparam signed [3:0] p15 = (-{((5'd30)|(-3'sd0)),(~&{1{(3'sd3)}})});
  localparam signed [4:0] p16 = {(-4'sd3),{1{{(4'd4)}}}};
  localparam signed [5:0] p17 = ((((5'sd14)&(3'd5))>=((-4'sd4)>>>(4'd3)))<=((6'd2 * (5'd6))!={(4'd5),(5'd21)}));

  assign y0 = ((p8?p15:p7)||(p10?p17:a4));
  assign y1 = ({4{$signed(p14)}});
  assign y2 = {3{((a4===a2)?(&a3):{3{a0}})}};
  assign y3 = {3{({2{p10}}+(+p2))}};
  assign y4 = {{{(|p9),(~|b0),(~^p10)},(~&(~&{(~|b3)}))}};
  assign y5 = (a0<<p11);
  assign y6 = (!{(3'd2),{{{p9}}},(4'd13)});
  assign y7 = (~(|{3{b3}}));
  assign y8 = (~($signed(((a5?a0:a1)|$unsigned((+(&p4)))))));
  assign y9 = (5'd6);
  assign y10 = (2'd3);
  assign y11 = ((~|((|(p12<<b5))>>>((~a5)>>>(p13!=p6))))>>((b5!==b3)*(p2<b4)));
  assign y12 = {((p0)),(~&$signed(b1))};
  assign y13 = {1{{3{({1{(2'sd1)}}^~{4{p4}})}}}};
  assign y14 = (p4<=p8);
  assign y15 = (-3'sd0);
  assign y16 = (!((a2===b0)>>>(-2'sd1)));
  assign y17 = (^($unsigned((-((~(b3==a1))>=(4'd11))))!==((-4'sd2)>((~|a1)!==(2'sd0)))));
endmodule
