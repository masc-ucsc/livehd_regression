module expression_00624(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-4'sd1)/(3'd5))>=(^((3'd6)?(-3'sd3):(4'sd7))))^((~((5'sd5)|(3'd5)))>>>(~^((4'd1)?(4'sd6):(4'sd0)))));
  localparam [4:0] p1 = {1{{(-3'sd3),(3'd5),(-3'sd1)}}};
  localparam [5:0] p2 = ({((&(-3'sd2))?(!(-2'sd0)):((2'sd0)?(5'sd9):(3'd7)))}>=((~|{(5'sd1),(3'd1),(3'd7)})<<((-4'sd4)^~(5'd21))));
  localparam signed [3:0] p3 = ((5'sd6)^~(2'd1));
  localparam signed [4:0] p4 = (6'd2 * ((4'd10)^(3'd1)));
  localparam signed [5:0] p5 = (((2'd3)^(4'd5))^~((-2'sd0)?(-5'sd8):(3'd3)));
  localparam [3:0] p6 = (-(((5'sd3)|(4'sd2))<((-5'sd0)+(5'd4))));
  localparam [4:0] p7 = (6'd2 * ((4'd13)==(5'd29)));
  localparam [5:0] p8 = (+(4'd15));
  localparam signed [3:0] p9 = (5'd4);
  localparam signed [4:0] p10 = (3'sd1);
  localparam signed [5:0] p11 = (3'sd1);
  localparam [3:0] p12 = ((5'd31)-((4'd9)===(-2'sd1)));
  localparam [4:0] p13 = {4{(-5'sd3)}};
  localparam [5:0] p14 = ((|(5'd25))==(-(((-4'sd7)<<(5'sd13))>((5'sd4)+(3'd1)))));
  localparam signed [3:0] p15 = (-3'sd1);
  localparam signed [4:0] p16 = {3{{3{(2'd0)}}}};
  localparam signed [5:0] p17 = (-3'sd2);

  assign y0 = {2{b0}};
  assign y1 = {1{((p1?a0:p1)?(p15?p6:p0):(^a5))}};
  assign y2 = (~(5'd27));
  assign y3 = {p15,p2};
  assign y4 = (5'd18);
  assign y5 = ({(a5?p13:a0)}>=(b4?a0:p14));
  assign y6 = {(p1^~a4),(^b0),(|a2)};
  assign y7 = (((p11>b4)?(a1>>>a3):($signed(p16))));
  assign y8 = $signed((~^(!(&a5))));
  assign y9 = (&((p2-p13)/a3));
  assign y10 = {p17,p7,p14};
  assign y11 = ($unsigned(((b4)&&(p17<=p16)))<$unsigned((5'd26)));
  assign y12 = (!{(5'd25),((a5===b1)>>{p0,p5}),{(~|p11),(b5^p17)}});
  assign y13 = (5'd20);
  assign y14 = (6'd2 * $unsigned((p15^~a4)));
  assign y15 = $signed({3{{2{{4{b3}}}}}});
  assign y16 = (-2'sd0);
  assign y17 = $unsigned($unsigned((~&(|(-(~|(-$unsigned({p6,p15,p0}))))))));
endmodule
