module expression_00947(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{{((5'd1)||(4'd9))}}};
  localparam [4:0] p1 = ((3'sd3)<<<(2'sd0));
  localparam [5:0] p2 = ((&({4{(-5'sd13)}}?(2'd1):(&(3'sd1))))!=={2{((-5'sd15)|(2'sd1))}});
  localparam signed [3:0] p3 = ((((2'd0)^~(2'sd0))-{(~^(3'd1))})>(!(~&(-((5'd15)?(2'd1):(4'sd3))))));
  localparam signed [4:0] p4 = (((2'd0)?(3'sd1):(2'sd0))?(&(5'd30)):(4'sd0));
  localparam signed [5:0] p5 = {{1{(!(!(-3'sd1)))}},{2{(!(2'sd0))}}};
  localparam [3:0] p6 = {2{({3{(5'sd3)}}^~((3'sd2)===(5'sd11)))}};
  localparam [4:0] p7 = (+((-2'sd1)?(3'd5):(2'd1)));
  localparam [5:0] p8 = (~^((((5'sd13)<<<(3'd2))?((4'd11)||(-3'sd1)):((2'd2)<=(3'd3)))^(((2'sd1)>=(5'd29))===((5'd14)?(5'd14):(-2'sd1)))));
  localparam signed [3:0] p9 = {3{(-{3{(5'sd10)}})}};
  localparam signed [4:0] p10 = {3{(((-3'sd2)&(5'd4))&((2'd2)>(4'd14)))}};
  localparam signed [5:0] p11 = (~(+(&(({(2'd2)}===(+(3'd0)))<({(2'd2),(3'd0)}===(~(-4'sd4)))))));
  localparam [3:0] p12 = (((+(5'd29))<<<((5'd29)^(3'sd0)))?((5'd18)?(-3'sd3):(5'sd9)):(((-2'sd0)?(5'sd15):(3'd6))-((3'd3)&&(4'sd1))));
  localparam [4:0] p13 = (~&((~|(~^(-((3'd4)^(-3'sd0)))))<<((+(2'sd0))>>>(^(2'sd1)))));
  localparam [5:0] p14 = (((3'sd2)<=(2'd0))^~(+((4'd1)?(4'd13):(-4'sd3))));
  localparam signed [3:0] p15 = (5'd29);
  localparam signed [4:0] p16 = (&(-2'sd1));
  localparam signed [5:0] p17 = ((+(4'd10))+(!((2'sd0)>=(5'd4))));

  assign y0 = $unsigned({p12,p4,p11});
  assign y1 = {(((a2<<b4)=={(b5?a2:p5)})|(~(4'd2 * {p7,b1})))};
  assign y2 = (~&(^(-4'sd5)));
  assign y3 = (+((|p9)!=(-p6)));
  assign y4 = {2{{3{p13}}}};
  assign y5 = {1{((~{2{{3{p10}}}}))}};
  assign y6 = (-({{p9,a2,a0},{p10,p11}}?(^(&(^(-p8)))):((-p9)?(p12?p8:p16):{p4,p9})));
  assign y7 = ((+(!(!p5)))<<((+p6)>>>{p4,p13}));
  assign y8 = (+(-{(!p1),(~^a2),(a0!==a3)}));
  assign y9 = (({a0}^(b2!=a4))?((a3^~a4)||(a2+b4)):((b0+a4)!==(b4==a3)));
  assign y10 = {4{(p12<=a1)}};
  assign y11 = {{4{b2}},((b5||b5)>>(a0>>>b4)),{(b4),(b3)}};
  assign y12 = ((6'd2 * (b2?a2:b0))?((4'd2 * b2)<=(b4||a2)):((~|a3)&&(b5<<b3)));
  assign y13 = (2'd1);
  assign y14 = (5'sd7);
  assign y15 = ($unsigned((+{2{(b0!==a1)}})));
  assign y16 = (~^((!((~^(~&b2))<=(&(b4+a1))))||(~((-(-b2))==((!p1))))));
  assign y17 = ((^((p5==b1)>>>(b2-p13)))-(-(&(p8<<p5))));
endmodule
