module expression_00628(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((3'd1)?(2'd0):(4'sd3)),{3{(5'sd5)}}};
  localparam [4:0] p1 = (&(((|((-5'sd9)+(5'sd13)))<<((2'd0)-(2'sd0)))&(((2'd1)==(4'd1))^((4'd0)>(-3'sd3)))));
  localparam [5:0] p2 = (-2'sd1);
  localparam signed [3:0] p3 = (-(|(((~|((2'd0)%(3'd2)))*((5'sd3)%(4'd2)))>>>(((-3'sd3)<<(-4'sd1))!=((3'd2)-(2'd3))))));
  localparam signed [4:0] p4 = (((5'd2 * (4'd11))>>((3'sd1)||(3'd4)))^~(((5'sd1)>>(5'sd15))&&((4'd10)<<<(2'd2))));
  localparam signed [5:0] p5 = (((4'd4)*(5'sd3))*((-3'sd3)!==(5'sd1)));
  localparam [3:0] p6 = (({(5'd15),(4'sd5),(-5'sd12)}<<((5'sd11)>>(-5'sd8)))<<<(((3'd2)==(-5'sd0))?(-4'sd5):((2'sd1)?(5'sd9):(2'sd0))));
  localparam [4:0] p7 = ((5'd2 * ((5'd29)?(4'd10):(4'd11)))-({(5'd12)}?((-4'sd3)||(5'd3)):{1{(5'sd5)}}));
  localparam [5:0] p8 = {((!((4'd1)!=(5'd25)))!={2{(+(-4'sd6))}}),({3{(4'd8)}}===(|(^{(5'sd12),(3'd7),(2'sd1)})))};
  localparam signed [3:0] p9 = ((!(4'd8))&&((2'sd1)?(-2'sd1):(5'd24)));
  localparam signed [4:0] p10 = (5'd29);
  localparam signed [5:0] p11 = (-4'sd5);
  localparam [3:0] p12 = ((4'd1)&(5'd10));
  localparam [4:0] p13 = (((4'sd4)?(-4'sd7):(4'd0))&((3'd2)<<<(2'd0)));
  localparam [5:0] p14 = (3'd7);
  localparam signed [3:0] p15 = (|(-{((3'd6)?(4'sd5):(2'd0))}));
  localparam signed [4:0] p16 = (~|{3{((4'd14)<(5'd18))}});
  localparam signed [5:0] p17 = {1{((5'sd11)?{3{(4'd3)}}:((-4'sd4)&&(5'd24)))}};

  assign y0 = {2{({4{b4}}!=(a0?p8:b1))}};
  assign y1 = (~&((&(!(^(~(a2==b2)))))?{(~|{2{b2}}),(b2>>b2)}:{4{(|a3)}}));
  assign y2 = (4'd3);
  assign y3 = $unsigned((-$unsigned((|$signed({2{a3}})))));
  assign y4 = ((-(~(-4'sd5)))^~((a5!=a4)!==(3'd3)));
  assign y5 = $unsigned($signed(b0));
  assign y6 = (3'd6);
  assign y7 = {{{2{$signed(b3)}},{(b5),{a0,b0,b4}}}};
  assign y8 = (2'sd0);
  assign y9 = {{(6'd2 * (b0<<b0))}};
  assign y10 = $unsigned($unsigned((|(~|(^(((|$unsigned((~&($signed((~|(~|$unsigned($unsigned($signed((^a0))))))))))))))))));
  assign y11 = ($signed({3{(-a5)}})>=$unsigned(((^$signed((b0<b2))))));
  assign y12 = {(2'd0),((p0==p5)>=(5'd19)),{((3'sd0)),{1{{p5}}}}};
  assign y13 = (a4?a5:a4);
  assign y14 = (!(((a0?b5:b2)?(4'd0):(a0?a5:b3))?(|(~(&(3'd1)))):((4'd3)?(b3?a0:a1):(a2?a0:b1))));
  assign y15 = (5'sd8);
  assign y16 = $signed(((~^(&(a5?b4:p14)))?(^$signed($unsigned((b5?b4:a2)))):($unsigned(a4)?(p7):(-a4))));
  assign y17 = (5'sd6);
endmodule
