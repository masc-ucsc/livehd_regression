module expression_00513(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'sd0);
  localparam [4:0] p1 = ((5'd30)==(6'd2 * ((3'd3)<<(5'd22))));
  localparam [5:0] p2 = {(((3'd0)?(3'd6):(-3'sd2))>>>(5'd2 * (4'd6)))};
  localparam signed [3:0] p3 = (({(2'd1)}&((4'sd1)?(3'd2):(-3'sd0)))<(3'd3));
  localparam signed [4:0] p4 = (-4'sd3);
  localparam signed [5:0] p5 = (4'sd0);
  localparam [3:0] p6 = (&((((3'sd3)?(2'd2):(4'sd0))||(!(5'd24)))?((-2'sd1)?(5'sd5):(5'sd4)):(2'd2)));
  localparam [4:0] p7 = (5'sd14);
  localparam [5:0] p8 = (~&(-(~^(~^(~^(5'sd9))))));
  localparam signed [3:0] p9 = {(5'd29),(-4'sd1),(5'd22)};
  localparam signed [4:0] p10 = (^(~|(~|((4'd12)!==(-5'sd14)))));
  localparam signed [5:0] p11 = (~|(((3'd5)||(2'd2))*(-4'sd5)));
  localparam [3:0] p12 = (-4'sd7);
  localparam [4:0] p13 = (!{3{{4{(-4'sd6)}}}});
  localparam [5:0] p14 = (+{2{((-4'sd3)==(3'sd1))}});
  localparam signed [3:0] p15 = ((&(5'd24))<=(~^(-5'sd6)));
  localparam signed [4:0] p16 = (-4'sd2);
  localparam signed [5:0] p17 = {4{{(2'd0),(4'd14),(2'd3)}}};

  assign y0 = $unsigned(($signed(((-(b3===a3))*$signed((5'd16))))));
  assign y1 = (~^{(+(~^((a5<p12)>(^a5)))),({{p9,b3}}>>(^{b1,p12,a1}))});
  assign y2 = (&(5'sd12));
  assign y3 = (&b1);
  assign y4 = {2{(~^(^(|a1)))}};
  assign y5 = (~^((b3<<<b2)>(|(!p13))));
  assign y6 = (2'd0);
  assign y7 = ((b4+a5)?(a3===b0):(~&(|b2)));
  assign y8 = ({{p6,p12,p10}}<<(p10?p12:p13));
  assign y9 = ((&(b0?a4:p5))<((p4!=p3)||{a3}));
  assign y10 = {1{(((b2?p5:p16)!={3{p3}})?(5'd2 * {3{b1}}):((p11?p16:p12)?{1{a5}}:(p11?p12:p9)))}};
  assign y11 = {3{((b2^~p6)&$signed((p7)))}};
  assign y12 = {((p10^p12)&{(b1|p4)}),({p2,p0,p2}^{1{(|a4)}}),{(~|(+(&(a1?a1:p5))))}};
  assign y13 = (((-(^b3))>>>(~(~a5)))?(-(~|$unsigned(((p8?p0:a1)|(b4>=b1))))):(~&((~|(a0?b3:p10))&&$signed((a0?p6:p10)))));
  assign y14 = (+(~(((p5?p11:p3)||{(p10^~a1)})<=((p4==p2)?(p17?p8:p17):$unsigned((p12))))));
  assign y15 = {(-(&(&{(~^({a3,b3,p6}?{{b3},(-a4)}:(|(a0?a5:p15))))})))};
  assign y16 = ((~&(~|(!(4'sd4))))?((&a1)?(|a3):(5'sd4)):((b5?a4:p4)?(b4?a0:b5):(a2+b0)));
  assign y17 = ((p4?p0:p10)*(p8));
endmodule
