module expression_00660(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(5'd28),(5'd7)};
  localparam [4:0] p1 = ({4{(5'sd12)}}?{3{(5'd8)}}:((5'sd14)?(2'sd1):(-3'sd0)));
  localparam [5:0] p2 = ((((4'd12)?(2'd2):(3'sd0))?((-5'sd7)?(4'd8):(5'd2)):((2'sd1)?(4'sd3):(4'd5)))?(((2'd0)?(-4'sd5):(2'd0))?((4'd2)?(3'd2):(4'sd3)):((4'd9)?(2'sd1):(-2'sd1))):(((-3'sd0)?(-4'sd1):(3'sd1))?((5'd30)?(-2'sd0):(-2'sd1)):((-5'sd13)?(3'd0):(3'd5))));
  localparam signed [3:0] p3 = (+((&{4{(2'd3)}})?{4{(3'd4)}}:(~&(-{1{(5'sd4)}}))));
  localparam signed [4:0] p4 = (!((&(-5'sd6))&&((-3'sd3)!==(2'd1))));
  localparam signed [5:0] p5 = (-3'sd3);
  localparam [3:0] p6 = ((((5'd18)!=(2'sd1))?((3'd3)?(5'sd3):(2'sd1)):(-2'sd0))&&((~|(2'd2))===((2'sd0)==(-4'sd2))));
  localparam [4:0] p7 = (4'd12);
  localparam [5:0] p8 = ((((2'd0)==(-4'sd5))>=((5'd3)?(4'd6):(4'sd5)))<<<(((-3'sd1)&(-3'sd3))>((5'd27)<<(2'sd1))));
  localparam signed [3:0] p9 = {4{(-4'sd2)}};
  localparam signed [4:0] p10 = (&(5'd18));
  localparam signed [5:0] p11 = ((((3'd7)!=(5'd5))*((3'd7)!=(3'd6)))-(|(~&(((-5'sd1)===(4'd13))!=(+(5'sd7))))));
  localparam [3:0] p12 = ((((2'd0)?(3'd1):(5'sd10))?((-3'sd1)?(3'd3):(3'sd3)):((-3'sd1)&&(2'd2)))!=((((3'd2)===(5'sd3))!=(&(2'sd1)))||({(5'sd1),(4'sd2),(2'd1)}-{(2'sd1),(5'd18),(2'd3)})));
  localparam [4:0] p13 = (|(~|(~^(-(~&(^(|(|(!(|(-(^(|(~^(~&(4'd6))))))))))))))));
  localparam [5:0] p14 = (4'd9);
  localparam signed [3:0] p15 = ((~&((4'd10)?(5'd16):(2'd1)))?((3'sd1)?(3'd2):(2'sd0)):((4'd7)?(-3'sd0):(4'sd3)));
  localparam signed [4:0] p16 = {1{{2{(5'sd11)}}}};
  localparam signed [5:0] p17 = {3{{3{(-2'sd1)}}}};

  assign y0 = ((4'd8)&(((~&p17)%b3)>>$unsigned((~|(p7!=a1)))));
  assign y1 = ({3{{1{p1}}}}|(-{(b3>=p4),(&b0),{2{a5}}}));
  assign y2 = ((&(a5?p9:b4)));
  assign y3 = (5'sd15);
  assign y4 = ((a2?p6:p10)?{(^b5)}:(a5?b1:p13));
  assign y5 = ((~^{2{(b1^~p13)}})&&((p9?p7:a3)&(+(b5?p11:a2))));
  assign y6 = ((-4'sd2)===((5'd2 * (5'd27))^~(b2?b3:b3)));
  assign y7 = {3{(5'd26)}};
  assign y8 = ((3'd5)^~((2'd0)|{4{p13}}));
  assign y9 = (~&{{{(p9>>p6),{p0,p16},{p13,p16,p12}}},({(4'd2 * p2),(p15>>>p10)}<<({p9,p1,p15}&&(p7|a2)))});
  assign y10 = ((p3&p13)>(p14>=p8));
  assign y11 = (5'd2 * (p8&a0));
  assign y12 = ((-2'sd0)&&(2'sd0));
  assign y13 = (-(~|(~|p4)));
  assign y14 = ({3{{b1,a4}}}==={(((a5&&b1)|{b1,b2,b0})!={2{$unsigned(b1)}})});
  assign y15 = $signed((~&{2{((|p13)?{4{p1}}:{p5})}}));
  assign y16 = {{{({4{p15}}^(-4'sd4))}},{{p14,p10},(p1+p3)},(-2'sd0)};
  assign y17 = ((p15?p15:p9)||(p11||p2));
endmodule
