module expression_00605(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(~|{1{{4{{3{(3'd1)}}}}}}));
  localparam [4:0] p1 = (~&(5'd27));
  localparam [5:0] p2 = (({3{(5'sd7)}}?((3'sd2)?(2'd1):(4'd9)):{2{(4'd4)}})-(6'd2 * ((2'd1)?(5'd3):(5'd31))));
  localparam signed [3:0] p3 = {1{{4{{1{{4{(3'sd2)}}}}}}}};
  localparam signed [4:0] p4 = (((2'sd0)?(4'sd3):(5'd18))?{(!((3'd5)?(5'd30):(2'sd1)))}:((2'd1)?(4'd6):(2'd0)));
  localparam signed [5:0] p5 = (!{(((5'sd10)>>(3'd2))>>>{(-3'sd1),(3'd4),(5'd20)})});
  localparam [3:0] p6 = ((((4'sd1)<=(-4'sd1))!=((-4'sd0)!==(5'sd2)))==(+{{(5'sd15),((5'd15)<=(5'd29))}}));
  localparam [4:0] p7 = {{2{(-3'sd1)}},{1{(3'd5)}},{3{(5'sd2)}}};
  localparam [5:0] p8 = (^{(3'd2),(3'sd3)});
  localparam signed [3:0] p9 = ({1{(~|((~{1{(-5'sd11)}})>>(+(+(5'd12)))))}}<=((((5'd17)+(2'd0))>(~|(4'd5)))>>>(~(+(~(3'd6))))));
  localparam signed [4:0] p10 = (5'd2 * ((4'd1)<<(2'd1)));
  localparam signed [5:0] p11 = (((-4'sd3)?(4'd5):(5'd31))?((3'd6)?(3'd7):(-4'sd3)):((2'd3)?(2'sd1):(5'd0)));
  localparam [3:0] p12 = (~^(~{(|{(-(2'sd1)),{(2'sd1),(2'd0),(3'd1)},{(2'd2)}}),((!(5'sd8))?((5'd3)?(2'd0):(-4'sd3)):{(5'd15)})}));
  localparam [4:0] p13 = (~^{4{{4{(-2'sd1)}}}});
  localparam [5:0] p14 = ((5'd2 * {4{(5'd27)}})-(((2'sd1)|(-4'sd1))?((5'd19)&&(2'd0)):{1{(2'd0)}}));
  localparam signed [3:0] p15 = ((((5'd22)>>>(4'd5))?((5'd22)===(4'd6)):(5'd2 * (3'd3)))-((3'd3)&&{3{(4'd4)}}));
  localparam signed [4:0] p16 = {((((5'd17)<<(-3'sd0))>=((2'd0)>(3'd0)))?(((-3'sd3)?(5'sd13):(2'd0))?(|(3'sd1)):{(-2'sd1),(3'd1)}):(~|({(4'd9),(-4'sd1),(4'd7)}<((4'd8)?(2'd2):(2'd2)))))};
  localparam signed [5:0] p17 = (^(5'd10));

  assign y0 = (~&(p10<=b2));
  assign y1 = ({(p12?a1:b2)}?$signed(({p11,p13}^$unsigned(a4))):((b3?p1:p16)>(p14&&p9)));
  assign y2 = ((p15?p12:p15)?(~&(p11?p7:b4)):(a2?p1:p7));
  assign y3 = {2{(-(-(~^{{2{p0}},(-p0),(~&b2)})))}};
  assign y4 = ((5'd8)^~{3{b4}});
  assign y5 = (((a1>>a1)===(b2^~a5))?{(p13?p4:a0),(a5?b0:a3),(a1===b0)}:((b0<p1)|(p7?p8:b1)));
  assign y6 = ({2{$signed(b1)}});
  assign y7 = (+a0);
  assign y8 = (&($signed({2{{3{p4}}}})+({3{p17}}==($signed(p17)<(p10>>p11)))));
  assign y9 = (({b4,p5}&(~$unsigned(p15)))!=$signed(((b2?p10:p15)?(+p10):{p5,p9,p12})));
  assign y10 = (&{1{{1{(~((p2?p3:b2)?(~p2):(~&p10)))}}}});
  assign y11 = $signed({3{(b4?p8:b5)}});
  assign y12 = {1{(((~&p9)?(p11<<<p14):(b1===b1))?{1{{{p15,p16,p5},(p15||a3),(p4>=p16)}}}:(~|{(a2?p3:p11),{p2},(&p11)}))}};
  assign y13 = (((~(a3<a0))?((a2===a1)<<(a0^a3)):$signed((b3/b5))));
  assign y14 = (6'd2 * {4{a2}});
  assign y15 = (-2'sd0);
  assign y16 = (+(^(^(p15<<<p17))));
  assign y17 = {4{(^p12)}};
endmodule
