module expression_00123(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+(3'd2))?{(5'sd2)}:(-4'sd1));
  localparam [4:0] p1 = (-((4'sd1)?(5'sd11):(-2'sd1)));
  localparam [5:0] p2 = ({((3'd3)?(-4'sd6):(5'sd7))}<=(((5'd24)?(4'd9):(-5'sd5))?((3'sd2)?(4'd10):(3'd4)):((4'd12)===(4'd14))));
  localparam signed [3:0] p3 = {1{((((3'd5)+(3'sd2))>>{1{((3'd4)^(5'd5))}})^((6'd2 * (4'd4))>>>{4{(4'sd1)}}))}};
  localparam signed [4:0] p4 = ((((2'd0)?(3'd7):(3'd5))!==(~^(4'd4)))?((3'd4)?(-5'sd15):(-5'sd8)):(~|((2'sd1)>>(4'sd6))));
  localparam signed [5:0] p5 = (-3'sd0);
  localparam [3:0] p6 = (&((((4'd4)*(3'd3))<((-2'sd1)>>(2'd1)))^~(((-4'sd0)?(2'd0):(-3'sd3))&&((2'sd0)==(4'd12)))));
  localparam [4:0] p7 = ((-(-{1{{4{(4'd12)}}}}))<={4{(-2'sd1)}});
  localparam [5:0] p8 = (!(|(&(4'd10))));
  localparam signed [3:0] p9 = (~(6'd2 * {{(3'd1),(4'd3),(4'd12)}}));
  localparam signed [4:0] p10 = (&(5'sd10));
  localparam signed [5:0] p11 = ((((2'd0)>>>(5'd12))<=(|(3'd2)))^(~^(((5'd21)<<<(5'sd1))<(-(-3'sd3)))));
  localparam [3:0] p12 = (((2'sd1)!=(5'sd2))*((-5'sd2)^~(5'sd15)));
  localparam [4:0] p13 = ((((-3'sd3)/(4'sd7))>((3'd1)%(2'sd0)))>>>((~((4'd10)===(5'd11)))/(-4'sd0)));
  localparam [5:0] p14 = {2{(-4'sd7)}};
  localparam signed [3:0] p15 = ((((-4'sd4)?(-4'sd0):(2'd3))==((3'd7)===(3'd5)))?((6'd2 * (2'd2))&&(4'd2 * (5'd30))):((3'd6)?(3'd0):(4'd9)));
  localparam signed [4:0] p16 = {1{{3{(5'sd12)}}}};
  localparam signed [5:0] p17 = (((~&((4'sd2)?(2'd0):(3'd7)))>>(^((5'd7)===(4'd2))))&{1{(((4'd13)&&(3'd7))>=(&(-5'sd4)))}});

  assign y0 = (~&(b2?a1:a0));
  assign y1 = {{(~&{p15,p3,a1}),{{a3},{p0,b3,b4}},(-(&{b3,a4,p0}))}};
  assign y2 = ($signed(a2)?(b1):(&a4));
  assign y3 = (~|((^(b0?p1:p6))>{1{(|(|p12))}}));
  assign y4 = (|(-(-(~&(~^p4)))));
  assign y5 = (((p3<=p8)?(b0!==b2):(p14?p2:p4))==((p7?p9:p5)?{2{p1}}:{3{p16}}));
  assign y6 = (^((^$unsigned((|(~|b4))))+(+{b2,p7,p15})));
  assign y7 = ({({p8,p15}<=(b1!==a1)),({p10,p14}>=(-3'sd3)),(3'd6)});
  assign y8 = (((p13<p12)&(p7>>>p14))<(~{{p5,p1,p12}}));
  assign y9 = ((b4?a1:b2)?(b3?a5:a5):(a4?b3:b3));
  assign y10 = (!{4{(a5)}});
  assign y11 = (p15>>p2);
  assign y12 = $signed((!(!(|(~|$signed(((a1^b2))))))));
  assign y13 = {(5'd4)};
  assign y14 = (|(p14<p12));
  assign y15 = ((^{1{((~^p3)>>>{p9,p2,p6})}})!=((p11|p11)<(+{p3,p8})));
  assign y16 = ((b2<<b0)+(a3?p1:b5));
  assign y17 = {{4{b0}},{3{b5}},(~|(b5?b0:b4))};
endmodule
