module expression_00603(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((!(!((^(2'd0))===((-2'sd0)<<(3'd6)))))==={1{((~|(3'sd2))>>(~|(-3'sd0)))}});
  localparam [4:0] p1 = {((-5'sd1)?(-2'sd1):(-4'sd1)),(|(-3'sd0)),{(3'd3)}};
  localparam [5:0] p2 = (((-5'sd8)>>>((3'sd3)===(-2'sd1)))<<<((5'd2)>>((-5'sd1)>=(-4'sd6))));
  localparam signed [3:0] p3 = (-5'sd4);
  localparam signed [4:0] p4 = ((((2'd0)>>(5'd13))!=((2'd2)|(-3'sd0)))<(((5'd14)?(3'd6):(2'd3))===((-2'sd0)^~(3'sd1))));
  localparam signed [5:0] p5 = (~|{2{(3'd4)}});
  localparam [3:0] p6 = ((2'd3)<<((2'd2)!==((5'd0)^~(-5'sd6))));
  localparam [4:0] p7 = ((-4'sd3)>(((3'sd0)>>>(3'sd2))||((3'd5)<<<(2'd1))));
  localparam [5:0] p8 = ((^((~|(5'd13))+((5'd7)>=(-2'sd1))))||{(&((-5'sd13)&&(-5'sd2)))});
  localparam signed [3:0] p9 = (2'd3);
  localparam signed [4:0] p10 = (({(5'd14)}&(+(3'd5)))?(!((2'd2)?(2'sd0):(5'd28))):{(5'd30),(3'd2),(2'd2)});
  localparam signed [5:0] p11 = (4'd10);
  localparam [3:0] p12 = (~|{((3'd6)!=(3'd5))});
  localparam [4:0] p13 = (^((~|(!((+(-2'sd0))>(~|(-3'sd3)))))>=(-(&(+(~^(^(2'd3))))))));
  localparam [5:0] p14 = (&(((5'd20)!=(3'sd1))&((3'sd3)!==(4'sd7))));
  localparam signed [3:0] p15 = (4'd2);
  localparam signed [4:0] p16 = ((((-5'sd4)<(3'd4))^~((5'd30)!==(-3'sd2)))^((+(5'd31))!=((3'd2)>>>(5'sd10))));
  localparam signed [5:0] p17 = (+(^((2'd2)?(2'd3):(4'd12))));

  assign y0 = ((((p15?p16:p17)!=(p8?a5:p15))==(a0?b2:p7))|{2{({1{p10}}>>>(p5<<p16))}});
  assign y1 = {(p12?b0:p4),(5'd2 * (4'd2 * b2)),(!((-3'sd2)))};
  assign y2 = (a5===a1);
  assign y3 = (|(-(-4'sd3)));
  assign y4 = (4'd12);
  assign y5 = (b0<<p5);
  assign y6 = (p10?p2:p5);
  assign y7 = (-4'sd7);
  assign y8 = {({p8,b3}^~{p7}),(5'd2 * (p7<p1))};
  assign y9 = {b4,a1,a2};
  assign y10 = {{{(2'd2)}},((b4||b4)-{b2,p6,a5}),(-3'sd0)};
  assign y11 = (((~|b4)?(p9?p15:b4):{p0})?((p10?p10:b3)!=(a0?p12:p13)):(~^({p3}?(~^p12):{p3})));
  assign y12 = $unsigned(((-4'sd4)));
  assign y13 = (5'sd1);
  assign y14 = (((!((&p16)>>{b2})))^~{(&b2),(b2|p8),$unsigned(p9)});
  assign y15 = {{(b2!==a5)}};
  assign y16 = {3{{1{(p10^~p16)}}}};
  assign y17 = (~(|($unsigned((~|{4{b3}}))<<(~^(b5>=a3)))));
endmodule
