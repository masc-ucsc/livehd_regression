module expression_00243(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({3{{(3'd1)}}}^~(~|({1{(5'd31)}}?((-3'sd2)?(4'd0):(-3'sd0)):((2'd1)<<<(3'sd0)))));
  localparam [4:0] p1 = (5'sd15);
  localparam [5:0] p2 = (~|(2'd1));
  localparam signed [3:0] p3 = (-3'sd0);
  localparam signed [4:0] p4 = (4'd14);
  localparam signed [5:0] p5 = (4'd13);
  localparam [3:0] p6 = (5'd2 * ((3'd4)||(3'd5)));
  localparam [4:0] p7 = {((2'd3)<(-5'sd14)),((2'd0)|(-5'sd10)),((5'd28)^(2'd3))};
  localparam [5:0] p8 = (3'd1);
  localparam signed [3:0] p9 = (~((~((4'd7)?(3'd4):(4'd11)))?((^(3'd3))*(~^(3'sd1))):(~|((5'd11)?(2'd3):(-3'sd2)))));
  localparam signed [4:0] p10 = (((4'sd6)^~(2'd0))|(-2'sd1));
  localparam signed [5:0] p11 = (~^(|({4{(|(3'd4))}}!=(-{{(4'd9),(2'd1)},((5'd13)&(2'd3)),((3'd4)?(3'd7):(-5'sd7))}))));
  localparam [3:0] p12 = ((((2'd3)?(4'sd7):(4'sd5))&&((-2'sd0)<<<(-3'sd1)))<((~(2'd0))>=((3'd1)?(3'd5):(4'sd7))));
  localparam [4:0] p13 = ((((3'd2)?(4'sd2):(5'sd13))?(^(5'd6)):(+(5'd6)))?(~^((2'sd1)?(5'sd6):(3'd5))):(((4'sd1)?(-3'sd1):(2'd1))?(~(3'd3)):(!(-2'sd1))));
  localparam [5:0] p14 = (~^((5'd3)<=(4'd11)));
  localparam signed [3:0] p15 = (~^(~^(~^{1{{3{{4{(4'd12)}}}}}})));
  localparam signed [4:0] p16 = {4{(-5'sd1)}};
  localparam signed [5:0] p17 = ((^(2'd2))^~((5'sd3)<=(4'd8)));

  assign y0 = (p5<<<p14);
  assign y1 = ((-{(a0<p5),(a2^b0),(~^b5)})<(&{(a3&&p8),(-p4),(p12+a5)}));
  assign y2 = {2{(&(~&$signed(a5)))}};
  assign y3 = $unsigned((({1{$unsigned((-2'sd0))}}!==(&{3{b2}}))>=({2{(5'd2 * b1)}}=={1{(a0<p11)}})));
  assign y4 = (|{4{({a1}-(~p13))}});
  assign y5 = ((+(3'd2))?(5'd25):(~(4'd9)));
  assign y6 = ((p15^a4)>>(b4<a1));
  assign y7 = ({(!(b5?p13:p6)),{(a2!==a3)},(p1^b5)}||({(p8<b5)}?(p15^a4):(a3-b5)));
  assign y8 = (($signed(((a4<<<b2)<<$signed(a2))))^(({4{b0}})-(a4&b2)));
  assign y9 = ($signed(({(p7&&p7)}&&($unsigned(p2)<<<$signed(p2))))>>>{{($signed({p14,p10})==({p14,p11,p7}))}});
  assign y10 = ((p15>b0)?(p7^p16):(p9?p2:p7));
  assign y11 = ($unsigned(((p3?p17:p9)%p5))<<<(4'd14));
  assign y12 = (~{p14,a5});
  assign y13 = (((-p0)^(|p16))^~{4{b2}});
  assign y14 = $unsigned((5'd15));
  assign y15 = ((5'd2 * {(b2||b2)})|(!{(-((b3<=p3)-(4'd2 * b1)))}));
  assign y16 = (((a0<<<p15)&{b3,a4})<<(6'd2 * (&(a1===b1))));
  assign y17 = (-3'sd2);
endmodule
