module expression_00086(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(3'd3)}};
  localparam [4:0] p1 = (~^(-(&(+(~|(-4'sd1))))));
  localparam [5:0] p2 = {((5'sd1)!=({(-2'sd0),(-5'sd9),(4'sd4)}>>(+(-5'sd15))))};
  localparam signed [3:0] p3 = (((-3'sd0)===(-2'sd0))>((3'd5)&&(4'sd4)));
  localparam signed [4:0] p4 = ((5'd13)?{4{(2'd0)}}:{2{(-4'sd2)}});
  localparam signed [5:0] p5 = ((((2'sd0)==(-3'sd2))<<{4{(4'd0)}})&({3{(4'sd5)}}>>((2'd1)||(2'd1))));
  localparam [3:0] p6 = ((3'sd1)?(2'd1):(-5'sd14));
  localparam [4:0] p7 = ((5'd13)<<<(5'sd9));
  localparam [5:0] p8 = ({2{(2'sd0)}}=={(2'd0),(2'd3),(3'sd1)});
  localparam signed [3:0] p9 = {3{{2{((5'd10)!==(4'd4))}}}};
  localparam signed [4:0] p10 = ((-3'sd0)?(2'd0):(5'd2));
  localparam signed [5:0] p11 = ((~(-5'sd7))<<<(-4'sd0));
  localparam [3:0] p12 = {1{(3'd3)}};
  localparam [4:0] p13 = (-4'sd7);
  localparam [5:0] p14 = {4{(4'd7)}};
  localparam signed [3:0] p15 = (+(-({(4'd0),(3'd1)}<((5'd18)<<<(5'd21)))));
  localparam signed [4:0] p16 = {3{((3'd0)-(4'd0))}};
  localparam signed [5:0] p17 = ((~|{(5'd29),(5'd6)})?(+(|(4'sd7))):{(4'd6),(-5'sd8),(-4'sd3)});

  assign y0 = (3'd3);
  assign y1 = {3{{4{{3{b2}}}}}};
  assign y2 = (+(!{a3,a3,a3}));
  assign y3 = ($unsigned(p4)<=(p15>>>p10));
  assign y4 = (~&((~^{1{((|(p7?b0:p10))<(^{1{b0}}))}})^{3{(!{4{a5}})}}));
  assign y5 = (((b3*b1)&(a1?a2:b4))&&(~^((a0?p11:p7)==(p8/b3))));
  assign y6 = (2'sd0);
  assign y7 = (3'sd3);
  assign y8 = ((-3'sd1)?(a2?a1:b5):(4'd6));
  assign y9 = ((({a5,a1,p6}^~(3'sd2))<<({p15,p1,p10}&{2{p1}}))^~(2'd0));
  assign y10 = (-2'sd0);
  assign y11 = ((~^(6'd2 * (a2!=p12)))!=(~^($signed(a2)!=={a0,b3})));
  assign y12 = (!(~^(~(~^(!((($signed(p10))?{3{a1}}:(p10<<p13))-((b5?a0:a3)?(&(a0)):{3{a4}})))))));
  assign y13 = ((((!a4)?(|a0):(~a5)))===((a0?a4:a4)-($signed((b1*b5)))));
  assign y14 = {$unsigned((!({a4,p1,p0}<(p12)))),({{(+p8)},(b5?p0:p10)})};
  assign y15 = $signed({3{p0}});
  assign y16 = ((b1&p15)?(6'd2 * a1):(b5?b2:p11));
  assign y17 = (((p11>>>p6)?{3{p12}}:{2{p5}})^((a5<<<p12)>=(p17==p6)));
endmodule
