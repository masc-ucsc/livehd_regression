module expression_00090(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(((2'sd0)*(5'sd7))*((4'd4)&&(4'd2))));
  localparam [4:0] p1 = {1{((((3'd3)!==(3'sd1))<=(~&(3'sd3)))^(((-5'sd0)|(3'sd2))!=((2'sd0)>=(2'd0))))}};
  localparam [5:0] p2 = (~&{4{{4{(2'sd1)}}}});
  localparam signed [3:0] p3 = {{(4'sd0),(4'd12),(4'sd2)},{{2{(-3'sd1)}},{3{(-4'sd6)}}},({(-4'sd0)}^~{3{(2'd1)}})};
  localparam signed [4:0] p4 = (~^((2'd2)+(~(((-2'sd1)<<(3'd4))<<(!(2'd3))))));
  localparam signed [5:0] p5 = ({4{(5'sd4)}}+({3{(2'd2)}}<<(4'd14)));
  localparam [3:0] p6 = (3'd2);
  localparam [4:0] p7 = {(~^(&(2'd2))),((3'sd1)?(2'd2):(4'sd0)),((4'sd2)===(4'd6))};
  localparam [5:0] p8 = ((4'd2 * {(3'd2),(2'd3)})^~((-(~&(3'sd1)))!={2{(3'd6)}}));
  localparam signed [3:0] p9 = (^(4'd8));
  localparam signed [4:0] p10 = ((-5'sd6)>>>(-3'sd3));
  localparam signed [5:0] p11 = (3'd0);
  localparam [3:0] p12 = {(-2'sd1),{3{(-4'sd6)}}};
  localparam [4:0] p13 = (-(((4'd2)?(3'd7):(2'd2))?(4'd3):(-((3'd1)?(3'd4):(3'sd1)))));
  localparam [5:0] p14 = {({(4'd9)}=={3{(5'd0)}}),(((4'sd1)+(-2'sd0))|((4'sd6)<<(3'd6))),{2{{1{(-4'sd6)}}}}};
  localparam signed [3:0] p15 = ((-3'sd0)&&(5'd26));
  localparam signed [4:0] p16 = (-({(-5'sd15)}<(+(2'sd0))));
  localparam signed [5:0] p17 = (&((~^(&{(2'd3),(-2'sd0)}))&&(((-4'sd2)!=(3'd1))>(~|(-2'sd0)))));

  assign y0 = (4'd1);
  assign y1 = (+(((p7^a4)>=(+p13))?((&a2)?(~&b1):(p1?a0:p11)):((^p6)?(b4===b1):(a0?p10:p9))));
  assign y2 = (2'd3);
  assign y3 = ((~&(5'd22))^(|(3'd4)));
  assign y4 = ({(-p8),(-b2),(2'd0)}<={{({3{b1}}==(4'sd3))}});
  assign y5 = ((p8?a4:p2)&&(|(p5?a4:p17)));
  assign y6 = (-5'sd10);
  assign y7 = ((~^({4{p6}}&&(~|(p0<<<p0))))?((p5<p13)?(p17+p10):(b2||a1)):((!(p0!=p7))-{1{(6'd2 * p2)}}));
  assign y8 = ({2{a1}}?(5'sd8):(a1?a4:a3));
  assign y9 = {({2{b3}}?(p16?b5:b2):(3'sd0))};
  assign y10 = {3{(3'sd0)}};
  assign y11 = (3'sd2);
  assign y12 = ({3{{p8,p7,b5}}});
  assign y13 = ($signed(({p12,a4}?$unsigned(a3):$unsigned(p7)))?(({a2,a4}?(b5?b5:a2):$unsigned(b4))):$unsigned(($signed(b2)?(a0?b5:a5):{b1,p1,b1})));
  assign y14 = (((&(a1?p4:p6))?(a2&&p14):(a4!==a4))!={({a1,p7,p1}||((b1==p7)>=(p6^b3)))});
  assign y15 = (((-3'sd1)<=(2'sd0))?($signed(b5)!=(a1?a3:p2)):(p4?a2:p12));
  assign y16 = {3{p11}};
  assign y17 = ((&(~^(~&(p6?p11:p4))))?(|(~(~|(p1?p3:p16)))):(^((&p17)?(+p17):(~^p17))));
endmodule
