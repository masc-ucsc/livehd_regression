module expression_00437(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd3);
  localparam [4:0] p1 = (~&(((4'd9)===(3'sd0))?((5'sd15)>(2'd0)):((-2'sd0)&&(-3'sd2))));
  localparam [5:0] p2 = ({3{(3'sd0)}}===((^(5'sd0))==((4'sd1)?(2'd0):(-4'sd6))));
  localparam signed [3:0] p3 = (~|(5'sd2));
  localparam signed [4:0] p4 = {2{(+{1{{(4'sd0),(3'sd0),(-4'sd1)}}})}};
  localparam signed [5:0] p5 = (~|(|(+(~((5'd8)>>(~((-2'sd0)!=(-5'sd4))))))));
  localparam [3:0] p6 = {2{(-3'sd1)}};
  localparam [4:0] p7 = (5'd21);
  localparam [5:0] p8 = ((3'sd3)?(-3'sd3):(-2'sd1));
  localparam signed [3:0] p9 = {4{{2{(-5'sd10)}}}};
  localparam signed [4:0] p10 = (((3'd6)&(-2'sd1))<{(3'sd0),(5'd8),(-5'sd12)});
  localparam signed [5:0] p11 = (((3'd6)===(3'sd3))?((4'd8)==(5'd5)):((4'sd0)?(4'd7):(5'd29)));
  localparam [3:0] p12 = {{(+(4'd10)),(^(3'd6))}};
  localparam [4:0] p13 = (!(3'sd0));
  localparam [5:0] p14 = {3{(((2'sd0)?(2'd1):(2'sd1))?((2'd0)|(3'd0)):((-3'sd0)<<(-5'sd8)))}};
  localparam signed [3:0] p15 = ({1{{(-3'sd1),(-3'sd0),(-4'sd6)}}}^~(4'sd6));
  localparam signed [4:0] p16 = (^(2'd2));
  localparam signed [5:0] p17 = (!(((3'd3)===(-2'sd0))+{3{(!(-3'sd0))}}));

  assign y0 = {4{a5}};
  assign y1 = ({(p15?p0:p8),(p14^~a0)}?(&{(a4?p3:p9)}):((p7?p2:p3)?(|p10):(b1?p15:p8)));
  assign y2 = (+(((-p5)?(|p14):(p0?p5:p12))>((p7?p10:p6)^~(p17?p1:p8))));
  assign y3 = (-4'sd4);
  assign y4 = {2{{3{p5}}}};
  assign y5 = (6'd2 * (~(p8^p0)));
  assign y6 = ((b1+a5)&&(~^b5));
  assign y7 = (|(~|((-{3{{4{p13}}}})-(|(|{2{(p10|p12)}})))));
  assign y8 = {$signed((~{3{{3{p17}}}})),{(~&{p7,b2,b3}),{4{p17}},{p10,a2}}};
  assign y9 = ((~^p15)?(p3&p3):(p2?p14:p0));
  assign y10 = (3'sd1);
  assign y11 = ((2'd0)?{(p2?b5:p12)}:((~p5)));
  assign y12 = (3'sd3);
  assign y13 = {((^(2'sd0))),{2{(p7?p3:p2)}}};
  assign y14 = (&(+{3{(|(~|(!(~a0))))}}));
  assign y15 = {3{p14}};
  assign y16 = ((a1===a1)?(a3|b3):(^p17));
  assign y17 = {(a3?b3:b1)};
endmodule
