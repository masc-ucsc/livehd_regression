module expression_00480(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~((~(((2'd2)+(-2'sd1))-((5'sd8)<<<(3'd4))))!=={(~(3'd6)),((4'sd7)<<(4'd9)),((2'd0)!==(-3'sd3))}));
  localparam [4:0] p1 = {3{((!(3'sd3))<={4{(-4'sd7)}})}};
  localparam [5:0] p2 = (((5'sd8)?(3'sd1):(4'd4))?(((-3'sd0)^(-3'sd0))%(4'sd4)):((5'd2)>>>((5'd11)?(4'd1):(4'd5))));
  localparam signed [3:0] p3 = (+(|{(4'd14),(3'd6)}));
  localparam signed [4:0] p4 = (({(3'd3),(5'sd1),(2'sd0)}<<<{2{(2'd2)}})>=((5'd25)?(5'd10):(3'd6)));
  localparam signed [5:0] p5 = ({(4'd2 * (4'd14))}==((-5'sd14)?((-5'sd8)>(3'd4)):(3'd6)));
  localparam [3:0] p6 = {1{{1{{2{((~|{3{(3'd6)}})<=(!((2'sd0)^~(-4'sd5))))}}}}}};
  localparam [4:0] p7 = (2'd3);
  localparam [5:0] p8 = ((5'd20)&((-4'sd2)?(4'd2):(-5'sd7)));
  localparam signed [3:0] p9 = {2{(5'sd0)}};
  localparam signed [4:0] p10 = {4{(2'd0)}};
  localparam signed [5:0] p11 = {1{(4'd2 * ((5'd8)>>(2'd3)))}};
  localparam [3:0] p12 = (~(((~^((2'd3)===(-5'sd5)))=={3{(5'd30)}})^~((~^((-2'sd1)!==(3'd5)))<<<((3'd7)>=(5'sd0)))));
  localparam [4:0] p13 = ((^{(3'd3),(5'd23)})&((5'sd10)<<(2'sd0)));
  localparam [5:0] p14 = ({3{((3'd5)>>(4'd6))}}?(((2'd2)<(4'sd1))!=((5'd16)^(-3'sd1))):({4{(4'd5)}}&&((2'd1)?(2'd0):(4'd12))));
  localparam signed [3:0] p15 = (2'd0);
  localparam signed [4:0] p16 = (5'd3);
  localparam signed [5:0] p17 = ((5'd30)-((-2'sd1)!=(|(4'sd0))));

  assign y0 = {{{p14,p1,p17},(p4|p6)},$signed($signed(((p8?p5:p10))))};
  assign y1 = (b2>=p0);
  assign y2 = ((!((b2===b0)<<<(b4?b5:b2)))>((a5|a1)<={2{b0}}));
  assign y3 = (({4{p1}})>=($signed(p10)<<(p17-b2)));
  assign y4 = {2{(^(3'd5))}};
  assign y5 = (~(~^(((~&(p1?p13:a0))<((p7>=p0)>=(!a3)))<((~&(a4?p7:p9))>>((+b1)>(!p5))))));
  assign y6 = {1{(p8?p0:p5)}};
  assign y7 = (5'sd8);
  assign y8 = (~^{$unsigned({$unsigned($unsigned((~|{b0,b0})))}),(-(^$unsigned(((|$signed((^a5)))))))});
  assign y9 = {4{p10}};
  assign y10 = (~^(~|(~&{2{{3{p6}}}})));
  assign y11 = (((b1?a4:b4)>>(4'd2 * a1))==={(b2&b3),(b2<<<b5)});
  assign y12 = ($signed(((3'sd0)?(a4|b2):(p4|a2)))?((3'd1)?(p8):(p2)):((5'd26)<<(5'd25)));
  assign y13 = ((b4^~b0)/p4);
  assign y14 = ((a5?a1:a5)!==(a3?b3:a3));
  assign y15 = (~|(~^(|{3{((p14<<b1)&(p17&&p17))}})));
  assign y16 = (~(+(a0^~a0)));
  assign y17 = (a1?a0:a0);
endmodule
