module expression_00065(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-4'sd1);
  localparam [4:0] p1 = (-(~&(^(~&(+(!(~&(&((~&(4'd4))<(+(4'd15)))))))))));
  localparam [5:0] p2 = ({(-3'sd2),(4'd3),(2'd2)}?(&(^(2'd3))):{(!(!(2'sd0)))});
  localparam signed [3:0] p3 = ((~^(|((3'd0)-{3{(4'd15)}})))<<<{2{(-2'sd0)}});
  localparam signed [4:0] p4 = (-((((5'd24)>(4'sd1))===((2'd0)&&(2'd2)))!==(((4'd2)?(5'sd15):(3'd5))-((4'd7)!=(-3'sd2)))));
  localparam signed [5:0] p5 = {1{{({(-3'sd1),(2'd0)}<=(~^{(-4'sd3)})),({3{(3'sd1)}}?((5'd9)&(5'sd14)):((-5'sd4)?(4'd9):(3'sd2)))}}};
  localparam [3:0] p6 = (((-4'sd1)?(4'sd6):(3'd3))^((2'sd0)+(5'sd0)));
  localparam [4:0] p7 = {(5'd25)};
  localparam [5:0] p8 = ((-2'sd0)?((2'd1)?(2'sd1):(-5'sd13)):((3'sd0)?(5'd0):(-5'sd6)));
  localparam signed [3:0] p9 = (+(3'd3));
  localparam signed [4:0] p10 = {(2'd1),(5'sd8),(-4'sd1)};
  localparam signed [5:0] p11 = {4{(~^{3{(3'd6)}})}};
  localparam [3:0] p12 = (4'sd7);
  localparam [4:0] p13 = ({3{(2'd2)}}?(|(!(~&(2'd3)))):((~&(4'd13))!==(|(3'd4))));
  localparam [5:0] p14 = (5'd2 * {(3'd6),(2'd1)});
  localparam signed [3:0] p15 = (2'sd1);
  localparam signed [4:0] p16 = {{(|(4'd0))},{2{(5'd20)}},{4{(2'd2)}}};
  localparam signed [5:0] p17 = {(2'd0),(3'sd3)};

  assign y0 = (~&$unsigned((~^((+$signed({3{b5}}))!=={4{{1{a1}}}}))));
  assign y1 = {1{a1}};
  assign y2 = ($unsigned(((b2?a1:a0)))!=((b4?b0:a0)?(5'd2 * a1):(a5?a1:a2)));
  assign y3 = ({{4{p14}},(2'sd1)}?(b3?b0:b1):((-4'sd1)<(a4!==a0)));
  assign y4 = {{({(a5<<<p7),(b1<=b2)}<{({b0,p14}|(p9>>b5))})}};
  assign y5 = ((p1>=b3)/b1);
  assign y6 = ((^((&b4)^{1{a1}}))?({p2,p9}^{2{p2}}):{((b1?b2:p14)>>>(b0!==a4))});
  assign y7 = (3'd5);
  assign y8 = ({2{p4}}|(p17>=b4));
  assign y9 = (&((6'd2 * (p6!=p0))>>{(p6&&p1)}));
  assign y10 = (+(~^(($unsigned((p3>p17))%p2))));
  assign y11 = ((4'd2));
  assign y12 = $signed($unsigned($signed($signed({4{$unsigned(b0)}}))));
  assign y13 = (~&(((5'd10))!=(4'sd6)));
  assign y14 = (((5'd0)));
  assign y15 = (((+(p7==p5))-({p16,p7,p12}>>>(p14+a5)))>>(5'd2 * (b0!==b1)));
  assign y16 = (((3'd0)!==(b4|a1))<<((p8<=p11)+(p15==a4)));
  assign y17 = (($signed((b4==p8))?(b0?p3:a1):$unsigned((-4'sd6))));
endmodule
