module expression_00230(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^(5'sd13));
  localparam [4:0] p1 = (5'sd13);
  localparam [5:0] p2 = (-5'sd13);
  localparam signed [3:0] p3 = (((|(!(4'sd1)))+{2{(3'd3)}})<<<(((-3'sd3)||(-4'sd3))+(&(~^(-3'sd1)))));
  localparam signed [4:0] p4 = ((^((-3'sd2)?(5'd6):(4'd2)))?((5'd27)?(2'd2):(4'd1)):(~|(~|(5'd14))));
  localparam signed [5:0] p5 = (-5'sd4);
  localparam [3:0] p6 = (((|(5'd8))?((2'd0)<<(3'd5)):((4'sd2)>>(-2'sd1)))&&(((-4'sd2)?(5'sd1):(5'd11))>=((-4'sd5)<<(-2'sd0))));
  localparam [4:0] p7 = (&(&(4'd7)));
  localparam [5:0] p8 = {(((5'd3)?(5'd14):(-3'sd2))?((5'd4)>>>(3'd7)):((-4'sd4)<(3'd2)))};
  localparam signed [3:0] p9 = ((3'sd2)!==(5'd19));
  localparam signed [4:0] p10 = (((6'd2 * (4'd11))>={1{((5'd15)<(5'd13))}})|(!((~^(+(4'sd1)))^~((2'sd0)+(5'd13)))));
  localparam signed [5:0] p11 = ((((2'd0)|(3'd1))<={3{(2'sd0)}})-{3{(6'd2 * (4'd2))}});
  localparam [3:0] p12 = {(((5'sd6)^(5'd21))?(3'sd0):(-4'sd4)),(~^(((4'd9)&(-5'sd13))<=(2'd2))),((~(2'd2))?((3'd1)!=(4'd10)):(3'd0))};
  localparam [4:0] p13 = {1{{4{((2'd2)?(-3'sd0):(-3'sd0))}}}};
  localparam [5:0] p14 = ({2{((4'd7)<(4'd4))}}&&((~(-3'sd3))!=(~^(-3'sd2))));
  localparam signed [3:0] p15 = (!((2'sd1)?(5'd16):(5'sd8)));
  localparam signed [4:0] p16 = (-3'sd0);
  localparam signed [5:0] p17 = (-(-((~(2'd1))?(^(5'sd15)):(~(4'sd1)))));

  assign y0 = ({3{(a4<=b4)}}-{(-p8),(p14^~b3),(p10>>>a4)});
  assign y1 = $signed($signed(((~&({3{$signed(p9)}}))>>>(+{({2{a5}}===(a4))}))));
  assign y2 = ($signed({2{$signed((b2^~p13))}})^{4{(b0<<<b5)}});
  assign y3 = ({{(2'd3)}}<<<(((5'd8)==={a1})<<(5'sd7)));
  assign y4 = ((^(b0?b1:a0))?((b4?p2:a1)==(b1)):{2{(b4?a4:b0)}});
  assign y5 = (($unsigned(((!a1)>>>(b0&&b4))))!==$unsigned(((-(3'd2))|(5'd6))));
  assign y6 = ((a3?p5:a5)-(2'd2));
  assign y7 = (^((b5>>>a3)?(b5?a4:a2):(a2==a3)));
  assign y8 = {2{(~^{{((-2'sd0)>{p1,b2,b5})}})}};
  assign y9 = ((p4&a5)>=(a1^~p7));
  assign y10 = {(((~^(b4||b3))^~(|(a1>>>a2)))-((b1-b3)===(~|{b3})))};
  assign y11 = {2{({1{(5'd10)}}===$signed((5'sd10)))}};
  assign y12 = ({4{(a0>=p12)}}^~{4{(b4==p9)}});
  assign y13 = ((~^(({2{p7}})+{3{p4}}))>>((~$unsigned((p14||a4)))^((b3!==b4)!=(|p13))));
  assign y14 = (((~(~|(|p16)))<{2{{4{p9}}}})<(^(~((b2-p2)&&(5'd24)))));
  assign y15 = {2{(-{1{(|(p5<p0))}})}};
  assign y16 = (((~^a4)?(&a5):{2{a0}})?{{3{b1}},(a1?a2:b0)}:{$signed($unsigned(a2)),$signed({4{b1}})});
  assign y17 = {b0,a2};
endmodule
