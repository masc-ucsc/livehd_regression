module expression_00317(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(2'd3),(2'd2),(4'sd2)},((5'd6)==(4'd14))};
  localparam [4:0] p1 = (|(|(-(^(|(~&(4'd8)))))));
  localparam [5:0] p2 = ({(~^(&(-3'sd3))),((3'sd2)==(3'd6))}<=(~&(((-5'sd1)?(2'd3):(4'd5))<<{3{(-4'sd1)}})));
  localparam signed [3:0] p3 = (~&((^((-2'sd0)?(-3'sd2):(5'd11)))?(|(|(5'd2 * (5'd6)))):((-(2'd1))>>((2'sd1)?(5'd6):(-4'sd2)))));
  localparam signed [4:0] p4 = {3{((-3'sd0)==(4'd0))}};
  localparam signed [5:0] p5 = (((~(-2'sd1))||(~&(2'd0)))<=((~(5'd1))^((5'sd11)===(-5'sd3))));
  localparam [3:0] p6 = (-(+(4'd2 * {1{(3'd2)}})));
  localparam [4:0] p7 = (({(2'd0),(3'd6),(5'd1)}?((5'd17)?(2'sd1):(2'd1)):{(3'd6),(-2'sd1),(4'd6)})?{((-2'sd1)<<(4'sd0)),{(-2'sd0),(5'd6),(3'd2)}}:({(4'd10),(4'd9),(4'd1)}-((3'sd2)^(5'sd1))));
  localparam [5:0] p8 = (((-5'sd9)?(-5'sd2):(3'd1))?((5'd14)<<(-3'sd2)):((3'd3)?(5'd7):(3'sd3)));
  localparam signed [3:0] p9 = (4'd5);
  localparam signed [4:0] p10 = (-3'sd1);
  localparam signed [5:0] p11 = ((^(&(^((^(5'sd13))*((2'd0)?(3'd2):(5'd4))))))<=(((-3'sd1)?(5'd27):(4'd0))%(3'sd2)));
  localparam [3:0] p12 = {2{(3'sd0)}};
  localparam [4:0] p13 = (4'd15);
  localparam [5:0] p14 = ({1{{(5'd12),(4'sd0),(5'd31)}}}^(((2'd1)|(5'sd4))?((3'sd0)^(2'sd0)):(!(2'd2))));
  localparam signed [3:0] p15 = (~(5'd2 * (+{2{(3'd0)}})));
  localparam signed [4:0] p16 = {(^{(-5'sd4),(5'sd8)}),(&((4'd11)===(3'sd2))),((3'sd2)>>>(2'd2))};
  localparam signed [5:0] p17 = ((3'd3)?(2'd2):(4'd13));

  assign y0 = ((((p17+p10)==(p9>p15))<((~p15)&(5'd2 * a1)))!=((!{(b1||a0)})===({a2}!==(^a5))));
  assign y1 = (~|(((b3<<<b0)?(b3*b0):(~b1))?(~|(b1?a3:p15)):(~&((~^b3)>>>(p8<b5)))));
  assign y2 = (+(^{3{(3'd0)}}));
  assign y3 = ((a2?b2:b1)?({a1,b3}=={a0,b3,b1}):{(b3?b0:b1)});
  assign y4 = ((!(~(b4?b0:a1)))&(&(~|(&(a3?a4:p3)))));
  assign y5 = ((~^(-p12))-(~^(+b0)));
  assign y6 = {$signed(a3),{a0,a1,b5},(5'd18)};
  assign y7 = ((3'd7)-{p0,p4});
  assign y8 = (a5?b3:b4);
  assign y9 = ((a5?a0:a1)?(^{b5,b4}):(~|(a2?b2:b4)));
  assign y10 = ((p11?p7:a1));
  assign y11 = (&(($unsigned(a5)%a2)>=((!b4)<=(p4||b2))));
  assign y12 = (&(({2{b2}}!==(~a5))));
  assign y13 = {4{(p11?p16:p7)}};
  assign y14 = ({4{{2{b1}}}}!==({3{b0}}>>>{3{a2}}));
  assign y15 = (^{3{a3}});
  assign y16 = (((~^b1)?(&a1):(4'd0))?(&(|(4'd13))):({b4}?(b2?a3:b0):(+a0)));
  assign y17 = {1{p6}};
endmodule
