module expression_00829(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^(({4{(3'd4)}}===(3'd5))>=(^{1{{2{(5'd13)}}}})));
  localparam [4:0] p1 = ({2{{3{(5'sd4)}}}}|(~&(-4'sd1)));
  localparam [5:0] p2 = {{{4{(5'd25)}},((4'sd4)==(-5'sd5)),{(3'd0)}},{(((-5'sd8)!==(5'sd5))>>((-3'sd3)<(5'sd15)))},{3{(~&(-5'sd4))}}};
  localparam signed [3:0] p3 = {(3'd5),((-2'sd1)-(5'sd0))};
  localparam signed [4:0] p4 = (~^(!(((-2'sd1)?(4'd9):(-5'sd14))?(((5'sd1)?(4'sd7):(2'd3))>>((-4'sd1)>(3'sd3))):(+(|((4'd6)?(3'd1):(3'd5)))))));
  localparam signed [5:0] p5 = (((5'd10)&(4'd0))?((3'd2)?(4'sd2):(3'd1)):((5'd13)<=(3'sd1)));
  localparam [3:0] p6 = (5'd2 * ((3'd0)?(2'd2):(4'd1)));
  localparam [4:0] p7 = {2{({{2{(4'sd6)}}}&((3'd4)<<(5'sd5)))}};
  localparam [5:0] p8 = (((-5'sd1)!=((-2'sd1)?(-3'sd3):(4'd7)))^~({(3'sd1),(5'sd14),(-2'sd0)}>>>(((2'd2)>>(-3'sd3))===(4'd2 * (5'd3)))));
  localparam signed [3:0] p9 = {4{(-5'sd2)}};
  localparam signed [4:0] p10 = (({3{(-4'sd5)}}?(~^(3'd2)):((2'sd1)>=(3'd0)))===(((-3'sd0)!==(-5'sd15))?{3{(-3'sd3)}}:{4{(3'd0)}}));
  localparam signed [5:0] p11 = ({2{(&{4{(2'd3)}})}}+(((3'd6)?(4'd10):(2'sd1))>>(2'd0)));
  localparam [3:0] p12 = (-4'sd2);
  localparam [4:0] p13 = {(5'd26),(-4'sd3),(5'sd3)};
  localparam [5:0] p14 = ((((2'd3)*(4'sd4))^((5'd9)/(-5'sd7)))<=(((-3'sd3)<(5'd14))==((5'd11)!==(5'd2))));
  localparam signed [3:0] p15 = ((2'sd0)-(2'd2));
  localparam signed [4:0] p16 = {{4{(5'd28)}},(~((-2'sd0)?(4'sd1):(5'd22)))};
  localparam signed [5:0] p17 = ({(4'd3),(4'd11),(-2'sd0)}&&(3'd5));

  assign y0 = $signed({(({(5'd2 * a0),(b4||p12)}||{p3,p14,p3})==($signed((a4&&p2))-((p4^~b5)|(a2>=b5))))});
  assign y1 = (-(((&$signed(p6))>=(p15<<p15))||((~&(b4^~a2))>>{(b5<<a3)})));
  assign y2 = ($signed(((2'sd0)?{1{(3'd4)}}:(a2?a3:a4)))&(2'd0));
  assign y3 = (-5'sd13);
  assign y4 = (!(2'd3));
  assign y5 = (~^{3{(-3'sd0)}});
  assign y6 = (((^(p0<<<p10))?(p12?p10:p2):(!(a3?p3:a3)))!={((~&p13)>=(p3?p7:p2)),((b5===b2)<(!p15))});
  assign y7 = (4'd1);
  assign y8 = (&((+(^p4))?(-(p1?p3:p6)):(p12?p4:p4)));
  assign y9 = ((((a4?a4:b5)&(b4?a2:a2))^~(-4'sd7))>(((-3'sd1)>>(b5===a2))>>>(3'd4)));
  assign y10 = (2'sd1);
  assign y11 = {{(^a5),$signed(a0),(b4)}};
  assign y12 = ((p15?a2:a4)+(^(~|(b4-a5))));
  assign y13 = ((((~a1)!=={a3,b3,b0})+({b3,a0}!=(a2>>>b3)))!=={((+a1)===(a3-a5)),((b1!==a4)>>$unsigned(a0))});
  assign y14 = ((b0<<b3)>(p3?p17:b3));
  assign y15 = (((p13>>>b5)<={3{a3}})?(p5?a3:b5):(a2?a2:a5));
  assign y16 = ((b1||a4)?(~(b0&b5)):(p4?a5:b3));
  assign y17 = {2{(({p15}>>{3{p3}})+{4{p7}})}};
endmodule
