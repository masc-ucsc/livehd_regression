module expression_00591(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({{(-3'sd1)}}==={(-3'sd3),(3'd1),(5'd7)})||(((3'sd3)&&(-3'sd1))<((4'd11)+(2'sd1))));
  localparam [4:0] p1 = (4'd2);
  localparam [5:0] p2 = ({1{((-4'sd3)?(2'sd1):(-5'sd6))}}?{1{{2{{4{(4'sd7)}}}}}}:(((2'sd1)?(2'd0):(2'sd0))?{2{(4'd6)}}:((4'd6)?(-3'sd0):(5'sd13))));
  localparam signed [3:0] p3 = {4{(-5'sd12)}};
  localparam signed [4:0] p4 = {4{(5'd7)}};
  localparam signed [5:0] p5 = (((3'd1)?(5'sd8):(2'sd1))<=((4'd2 * (2'd2))===((2'sd1)<(-5'sd5))));
  localparam [3:0] p6 = ((-2'sd0)>>>((5'd2 * (2'd0))-((2'd1)>>(5'sd5))));
  localparam [4:0] p7 = {((5'd2 * ((3'd6)||(5'd8)))>>>(&{(+(2'sd0)),(+(4'd7)),(|(2'd1))}))};
  localparam [5:0] p8 = (((&{(-4'sd5),(5'sd8),(-5'sd3)})<=((4'd8)&&(2'd1)))||{{(5'd25),(5'd6),(5'd12)},(+{(4'sd1),(-3'sd1),(5'sd10)})});
  localparam signed [3:0] p9 = (5'd20);
  localparam signed [4:0] p10 = (+{((-5'sd12)?(-4'sd5):(2'd3)),((4'd6)<<(5'd17))});
  localparam signed [5:0] p11 = (2'd0);
  localparam [3:0] p12 = {{((|(~&(3'sd0)))<<((3'd7)>>(2'd2))),(~^(~{((5'd6)^~(4'd0)),(|(3'd6))}))}};
  localparam [4:0] p13 = ((+{1{(-4'sd4)}})?{1{(3'd5)}}:{1{(+(4'sd6))}});
  localparam [5:0] p14 = (2'sd1);
  localparam signed [3:0] p15 = (2'd3);
  localparam signed [4:0] p16 = (({(-2'sd1),(3'd4),(4'd8)}-{((5'sd10)&(4'd11))})^(((5'd19)^(5'sd4))?((4'sd6)?(3'd0):(3'sd1)):((-5'sd15)?(2'd1):(3'sd3))));
  localparam signed [5:0] p17 = (5'd5);

  assign y0 = {{(~&b4)},{3{p8}}};
  assign y1 = (((p6>b0)?(p14+p8):(p2?p9:p8))!=((p3?p12:p9)>=(~(!(~|p2)))));
  assign y2 = (((b0===b2)>=(b0|b1))!==((b0-b3)-(a2>=b1)));
  assign y3 = (((2'sd0)?(p12?b2:p8):(p15))?((~^(p9|p16))|((p1&&p0))):(5'd21));
  assign y4 = (^(3'sd0));
  assign y5 = (3'sd2);
  assign y6 = ($signed((-a4))?(&$unsigned(a3)):(p10>b0));
  assign y7 = (p11>=p17);
  assign y8 = {{((2'sd0)<(3'd0)),((a5>>>b5)===(b1<=a2)),(!(4'd5))}};
  assign y9 = (((+a4)-(a1>=a0))?(~^(a1&&a3)):(5'd2 * (a0?p13:b2)));
  assign y10 = (&(~^(&((~^((|(b1<=a2))>>(a1|a4)))^(&(!((a2^b4)|(~&(^b0)))))))));
  assign y11 = (~{4{b4}});
  assign y12 = (!(p6?b4:b0));
  assign y13 = {3{(4'd15)}};
  assign y14 = ((~^(~^b3))>>(b1+p1));
  assign y15 = {2{((~&a3)?(^a0):(5'sd13))}};
  assign y16 = {{4{((a1&&a2)<(p6?b4:b3))}}};
  assign y17 = (~&(5'sd11));
endmodule
