module expression_00511(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd3)>>(3'd4))>=((5'd2)>=(4'd10)))?(~&(~|((-4'sd5)?(3'sd3):(3'd7)))):(^(^(~^((3'd5)<=(2'd1))))));
  localparam [4:0] p1 = (((3'sd1)&&((2'sd1)==(-5'sd13)))-((5'd2 * (3'd5))<<((4'sd1)/(-3'sd1))));
  localparam [5:0] p2 = ((4'd5)>>((-4'sd6)?(5'd25):(3'd5)));
  localparam signed [3:0] p3 = {1{((((5'd31)?(4'sd7):(-5'sd10))?((3'sd3)===(3'sd2)):(3'd5))!=={2{{2{(3'sd2)}}}})}};
  localparam signed [4:0] p4 = {((-4'sd5)+(5'd19)),((-5'sd4)?(2'd0):(4'd5)),((2'd2)?(5'sd6):(3'd2))};
  localparam signed [5:0] p5 = (!(+(^((3'd6)>>((^(2'd3))^~((5'sd6)&&(3'sd1)))))));
  localparam [3:0] p6 = (4'd11);
  localparam [4:0] p7 = ((((2'sd1)?(5'd25):(5'd4))>=((-4'sd4)%(-5'sd3)))?(((3'd4)===(3'd1))?((3'd4)?(4'd12):(5'd28)):((-5'sd4)>>>(-4'sd5))):(((5'sd5)?(5'sd11):(2'd0))?((-2'sd1)<(2'sd1)):((3'sd3)?(4'sd3):(-5'sd14))));
  localparam [5:0] p8 = {3{{(5'd25),(-4'sd2),(5'd0)}}};
  localparam signed [3:0] p9 = ((((5'sd9)?(3'd4):(-4'sd6))!==((2'sd1)===(4'd8)))<=(((3'd6)^(2'd3))&&(+{(-2'sd0),(2'd0)})));
  localparam signed [4:0] p10 = (5'sd0);
  localparam signed [5:0] p11 = (2'd0);
  localparam [3:0] p12 = ((4'd2 * {(4'd2),(3'd0),(4'd6)})?((2'd2)?{(2'd3)}:((3'd3)<<(2'sd1))):(+{(2'sd1),(5'd22),(4'd7)}));
  localparam [4:0] p13 = (((~^((5'sd11)/(2'd3)))<<<(~|(!(4'sd7))))^~((&(+(4'sd2)))^~(~&((5'sd12)<<<(4'd6)))));
  localparam [5:0] p14 = (+(~&({((~&(~^(5'd31)))===((5'd26)!=(2'sd0)))}<<(|((~^(-(5'd20)))>={((5'd11)|(-2'sd0))})))));
  localparam signed [3:0] p15 = (~|(({3{(2'd0)}}<<<{1{(5'sd7)}})&&({3{(2'sd0)}}>=((4'sd3)|(4'd3)))));
  localparam signed [4:0] p16 = (3'd3);
  localparam signed [5:0] p17 = (((~&(2'sd1))<=(~&(3'd3)))^~((4'd2 * (3'd5))>((3'sd2)===(2'sd1))));

  assign y0 = (((p6?p1:p7)&(p10?p11:p0))?{((5'd20)?(p5>>p16):(p15+p10))}:((p0?p7:p3)<<(b3!==b0)));
  assign y1 = (-2'sd1);
  assign y2 = {({a1,b1}+(b4^~p6)),((a1!=p2)<<(a1>>a5)),{((a3>>a2)>>>(a4<<b4))}};
  assign y3 = (((~b5)>>(b4&&b1))>>((b1<<b0)>{b4,b5,a3}));
  assign y4 = (~{1{((~&(~&((|(-{1{(~&{3{{1{p17}}}})}}))))))}});
  assign y5 = ((!$unsigned((((4'd2 * p1)?(-b0):(~^a3)))))>>(({4{a0}}>(~p16))>>>{3{(a2!==b3)}}));
  assign y6 = (p15?p6:p6);
  assign y7 = {{p3,p9,p12}};
  assign y8 = (($signed(b2)||{4{a5}})?((b5?a3:b3)^$signed(b2)):((b4)==(p4>b3)));
  assign y9 = (~|($signed(((a1!==b0)*(p5<=p11)))!=($unsigned((p5*b2))?(p3>=p13):$signed((b4)))));
  assign y10 = (4'd12);
  assign y11 = (((2'sd0)!==(4'd0))||((a0^~p3)?(-2'sd1):(p10%p0)));
  assign y12 = (^(^(&(~|(4'sd1)))));
  assign y13 = (~^((^$unsigned((b5+a0)))<=(~&(p16^~p6))));
  assign y14 = $unsigned((((a1&&b0)&&(b2==b1))|{{b4,b2},(a4?b2:b0)}));
  assign y15 = (4'd1);
  assign y16 = {{b2,b0,a0},(|(^{b4,a5,a5}))};
  assign y17 = {4{{3{p1}}}};
endmodule
