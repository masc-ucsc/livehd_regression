module expression_00600(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{({2{(5'sd14)}}<<((5'd20)?(3'd1):(4'd13)))}};
  localparam [4:0] p1 = {{(((2'd3)==(3'sd0))>=((3'd2)?(4'sd3):(2'd3))),{((-4'sd2)?(2'd0):(2'd2)),{(2'd2),(4'd13)}}}};
  localparam [5:0] p2 = (4'sd6);
  localparam signed [3:0] p3 = {((4'd10)&&(2'd1)),((3'd2)?(5'sd0):(5'sd0)),((5'd27)!==(-4'sd6))};
  localparam signed [4:0] p4 = ((((4'sd1)===(-5'sd0))||((-5'sd1)?(3'sd0):(-3'sd0)))?(((3'sd3)?(-4'sd6):(3'sd2))!=((5'd31)?(5'd17):(-2'sd0))):(((-3'sd2)+(2'd0))^((3'd6)>(-2'sd0))));
  localparam signed [5:0] p5 = {((-5'sd14)?(5'd26):(2'd2)),(^(2'd0))};
  localparam [3:0] p6 = {((5'sd11)!==(-2'sd0)),((4'd2)>=(5'd22)),(~(3'sd1))};
  localparam [4:0] p7 = (((|(4'd0))?(4'sd2):{(2'sd0),(3'd2)})?(4'sd1):({(4'd4),(4'd2),(-4'sd1)}!==((5'd13)==(-4'sd4))));
  localparam [5:0] p8 = {1{(((5'd7)?(-5'sd11):(2'd3))?((-5'sd13)?(-3'sd1):(2'd3)):((5'd25)?(5'd30):(5'd0)))}};
  localparam signed [3:0] p9 = (((^((4'sd5)?(4'd15):(2'sd0)))|((5'd20)?(5'd8):(5'sd10)))<<((+(~^(-4'sd7)))||((-2'sd0)<<<(4'd1))));
  localparam signed [4:0] p10 = (~(+(((3'sd3)+(-3'sd0))*(^(!(4'sd7))))));
  localparam signed [5:0] p11 = (~(2'd2));
  localparam [3:0] p12 = {1{((((-3'sd0)|(4'd2))?(4'd4):(5'sd0))-(((-5'sd6)||(3'sd0))?((-3'sd2)^(-4'sd0)):((-2'sd0)?(2'd1):(4'd12))))}};
  localparam [4:0] p13 = (((2'd1)==(^(3'd6)))<=((!(4'sd6))!=(~|(3'sd3))));
  localparam [5:0] p14 = {(((5'd1)&(4'sd6))?(|(5'd11)):(!(4'd1)))};
  localparam signed [3:0] p15 = (~|(~|{(3'd5),(2'd2),(-3'sd0)}));
  localparam signed [4:0] p16 = (4'd9);
  localparam signed [5:0] p17 = ((5'd25)<<(4'd11));

  assign y0 = (((+((~|p2)*(&p15)))^~((p16==p4)<<<(p6!=p4)))+(6'd2 * (a2^b2)));
  assign y1 = ((6'd2 * a1)^~(~&{2{a4}}));
  assign y2 = ((b1||p14)^{a1});
  assign y3 = (p2<<<p5);
  assign y4 = (-({4{p4}}?(~&{2{(p10?p16:p15)}}):((p8?p11:p3)?(|p16):(~^p13))));
  assign y5 = {1{(6'd2 * (p13>>>p0))}};
  assign y6 = (+(2'sd0));
  assign y7 = (p3?p11:p2);
  assign y8 = (!((~&$unsigned((3'd4)))<<<(($unsigned($unsigned((^(+p10))))))));
  assign y9 = (3'd5);
  assign y10 = (((+(!(p0>p8)))^({4{b0}}||(b1^p14)))<<<(&{4{(a5^~b0)}}));
  assign y11 = {4{(b1==a5)}};
  assign y12 = {2{(~&a3)}};
  assign y13 = {4{b5}};
  assign y14 = (4'd9);
  assign y15 = (4'sd6);
  assign y16 = (3'd4);
  assign y17 = ({p13,p0}-(a2!==b1));
endmodule
