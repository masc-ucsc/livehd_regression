module expression_00822(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{((-2'sd1)?(-2'sd0):(3'd1))}};
  localparam [4:0] p1 = {(+(&(((+(-4'sd7))>>>((4'd10)>>>(-4'sd7)))<<(&({(4'd4),(3'sd2),(5'd2)}!=((-2'sd0)<<(5'sd14)))))))};
  localparam [5:0] p2 = ((~((+(3'd6))^~(&(5'sd9))))>(~^((~^(5'd14))?(~&(3'd5)):((2'd2)||(5'd21)))));
  localparam signed [3:0] p3 = (~&(-2'sd1));
  localparam signed [4:0] p4 = {4{(2'd2)}};
  localparam signed [5:0] p5 = (5'd2 * ((5'd5)-(2'd2)));
  localparam [3:0] p6 = (((-3'sd2)&&(5'sd3))<(~&(5'd6)));
  localparam [4:0] p7 = ((((2'd1)?(5'd3):(3'd5))>>((5'sd5)?(2'sd1):(4'd11)))<<<({2{(3'd3)}}>>(~|(~(-4'sd4)))));
  localparam [5:0] p8 = ((((-2'sd1)<<<(3'd0))!={2{(2'd3)}})||((-3'sd2)^~((3'd2)==(-3'sd2))));
  localparam signed [3:0] p9 = (-5'sd12);
  localparam signed [4:0] p10 = {4{((4'd10)^~(-2'sd0))}};
  localparam signed [5:0] p11 = ({(4'd14),(3'd5),(-3'sd3)}==({(3'd2),(5'sd3),(2'd3)}&((3'sd1)&(3'sd2))));
  localparam [3:0] p12 = {2{((4'd6)?(4'sd4):(3'd3))}};
  localparam [4:0] p13 = ((-3'sd2)?(3'd2):(5'd26));
  localparam [5:0] p14 = (2'd0);
  localparam signed [3:0] p15 = (+(~^{{(5'sd14),(-2'sd0),(-4'sd7)},{(2'sd0)}}));
  localparam signed [4:0] p16 = ((^(~((5'd29)?(4'd10):(3'sd0))))?(~^(~^(3'd2))):(3'd7));
  localparam signed [5:0] p17 = ((5'sd3)?(2'sd1):(2'sd1));

  assign y0 = {{2{a4}}};
  assign y1 = (((a0?b5:b2)>>(3'd4))?(-5'sd8):{{a1,p15},(2'd3),(b1<<p10)});
  assign y2 = (2'sd0);
  assign y3 = ((+p1)?{1{p3}}:(&p15));
  assign y4 = ((((&p10)||{p13})||{(3'd7),(+p11)})^(~|{$unsigned((3'sd2)),((p5<<p6)+(p15))}));
  assign y5 = ({(p6==p9),{p4,p12}}|((p9>b2)>=(^p2)));
  assign y6 = {{(b5>>>a4),(|{a1,a1})},((|(~&b1))^~(a5===a4))};
  assign y7 = (4'd0);
  assign y8 = ({((-3'sd2)>((-a3)^(!a4)))}<<<({p9,a3,a3}>=$unsigned((p16>>a5))));
  assign y9 = (((p16-a2)?{3{b2}}:(b4^~a1))>((a5^~p9)>>{1{b4}}));
  assign y10 = (4'd8);
  assign y11 = (~^(~&(!{(~&(^((~&p13)<(p16?b1:p15)))),((~|(b0?b0:a5))===(a4?a4:a2)),(|((p2?p15:a3)^(a5?b3:p12)))})));
  assign y12 = ((a0%b4)&&(p17<<a0));
  assign y13 = (~(&(~{((~&(|(!(5'd13))))?(2'sd1):{(|p5),(-p17)})})));
  assign y14 = (|(-(4'd2 * (p8==a0))));
  assign y15 = (2'sd1);
  assign y16 = (|(^(~(~^(+(|(~&(~(!(~&(+(~(|(-(~|(+(~|(-p2))))))))))))))))));
  assign y17 = ((b2?p13:a3)<<{1{(^a1)}});
endmodule
