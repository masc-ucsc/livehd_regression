module expression_00381(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd3);
  localparam [4:0] p1 = {(4'sd4),(3'sd1)};
  localparam [5:0] p2 = {{(3'd2),(4'd8),(3'sd3)},(5'sd14),{(2'd2)}};
  localparam signed [3:0] p3 = (4'd9);
  localparam signed [4:0] p4 = (((4'sd5)&(-2'sd0))?((4'sd6)&(4'sd7)):(~&((4'd6)>=(2'd3))));
  localparam signed [5:0] p5 = (^(5'sd9));
  localparam [3:0] p6 = ((((5'd19)<(3'd7))>=((4'd3)>>>(2'd1)))&&({(4'd12),(-2'sd0)}>=((4'sd0)+(2'd0))));
  localparam [4:0] p7 = (~(^(|(|(((5'd26)?(4'sd2):(-2'sd1))?((5'sd7)?(2'sd0):(-3'sd0)):(&(~^(-2'sd0))))))));
  localparam [5:0] p8 = {1{({1{((4'd12)<=(2'd1))}}?{(^(5'd24)),((-5'sd2)!==(5'sd2))}:((2'd0)?(-5'sd10):(-3'sd0)))}};
  localparam signed [3:0] p9 = (4'sd7);
  localparam signed [4:0] p10 = ((4'd8)!=(~|(^(2'd2))));
  localparam signed [5:0] p11 = {(6'd2 * ((2'd0)+(2'd2)))};
  localparam [3:0] p12 = {({{(-5'sd0),(3'd6),(2'sd1)}}<<(~^{(4'sd3)})),(+(5'd2 * {(4'd4),(4'd13),(3'd0)}))};
  localparam [4:0] p13 = ((|((2'sd0)?(4'sd2):(2'd3)))==(((4'd4)?(4'd4):(5'sd8))<={(2'd3),(2'd0),(-4'sd7)}));
  localparam [5:0] p14 = ((((2'sd0)>>>(3'd3))>>>{((2'd0)?(5'd7):(4'd10))})|(((-4'sd5)===(-3'sd2))>>((4'd6)?(-2'sd0):(3'd2))));
  localparam signed [3:0] p15 = {3{(4'd2 * (4'd1))}};
  localparam signed [4:0] p16 = ((|(3'sd3))?((4'sd3)?(3'sd2):(2'd2)):(~^(4'sd1)));
  localparam signed [5:0] p17 = ((-4'sd5)||(4'sd7));

  assign y0 = (({1{p14}}>={1{p2}})>(^{3{b0}}));
  assign y1 = (^({b1,b2,b2}?(p16?b2:a4):(a4||b0)));
  assign y2 = {4{(b5&&p4)}};
  assign y3 = $signed($unsigned($signed($signed($unsigned(($signed(($signed($signed(($signed($unsigned($signed($unsigned($signed($signed((($unsigned(a1))))))))))))))))))));
  assign y4 = (((-p12)&&(p10&&p11))>>((a3?a1:a5)===(b3==b0)));
  assign y5 = (a5&p5);
  assign y6 = {1{{3{(a5+b2)}}}};
  assign y7 = (3'sd3);
  assign y8 = {((a2<a4)==(6'd2 * a2)),{(a0<=b3),(b0|b5),(a4&a1)},({b2,a0,a0}>={a4,a4})};
  assign y9 = {2{{4{b4}}}};
  assign y10 = (^p4);
  assign y11 = {{{(2'sd1)},(a5^b3),(p3<<<a0)},((3'sd1)>>>(2'd3))};
  assign y12 = {$unsigned($unsigned($unsigned((($unsigned((b0>b3))||(b4<<<p14))^~{(4'sd1)}))))};
  assign y13 = (~^(((&$signed((~^{1{(p2)}}))))<<((~&{4{p0}}))));
  assign y14 = {(3'd1),((p13>>p12)||(~(p12+p14)))};
  assign y15 = {1{({(b1<=p2),(b0?a4:p7)}&&{2{(p1|p10)}})}};
  assign y16 = (&((-$signed((-(b4?a1:a1))))&((6'd2 * b2)===(a4?a4:a0))));
  assign y17 = ({2{{3{p2}}}}>>{1{($signed((p9==p3))<<<$signed({(a5<=p4)}))}});
endmodule
