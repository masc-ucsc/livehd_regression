module expression_00807(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd7);
  localparam [4:0] p1 = ({1{{(5'sd12),(5'd18),(3'd7)}}}!=={{3{(2'd3)}}});
  localparam [5:0] p2 = {(5'd8),(3'd5)};
  localparam signed [3:0] p3 = (~((-4'sd6)>=(4'sd6)));
  localparam signed [4:0] p4 = (({4{(2'd0)}}+(-{2{(4'd12)}}))+(|((|{3{(5'sd14)}})<<(~|((2'd3)>>>(-2'sd1))))));
  localparam signed [5:0] p5 = {(4'd14),((2'sd1)-(2'd3)),{(4'sd1),(3'd0)}};
  localparam [3:0] p6 = {3{(-2'sd0)}};
  localparam [4:0] p7 = (3'd1);
  localparam [5:0] p8 = (5'd21);
  localparam signed [3:0] p9 = (3'sd3);
  localparam signed [4:0] p10 = ((((3'sd1)/(3'd1))>=((4'd14)?(5'd21):(3'd1)))!=(4'd2 * ((5'd5)<<<(4'd12))));
  localparam signed [5:0] p11 = ({1{{(5'd25),(-4'sd7),(3'd0)}}}&&(&(((3'd4)?(2'sd0):(2'd3))||(4'sd6))));
  localparam [3:0] p12 = ({1{(~^({3{(3'd7)}}?(&(2'd1)):((2'd0)&(-2'sd0))))}}&{(((2'd2)&&(-5'sd13))^~((3'd3)?(5'd5):(2'd0)))});
  localparam [4:0] p13 = ((4'd2 * (4'd9))<((4'sd1)&(5'd0)));
  localparam [5:0] p14 = (((3'd1)<<<(5'd4))?(3'sd2):(2'd3));
  localparam signed [3:0] p15 = (^(2'd1));
  localparam signed [4:0] p16 = (~|{{(2'd1)},((2'sd1)?(4'd11):(5'd29)),{1{(-2'sd0)}}});
  localparam signed [5:0] p17 = (~&(({(3'sd2)}<<<(2'd0))!=((5'd29)?(-2'sd0):(3'sd1))));

  assign y0 = {1{((|((a4>b3)?(b1?a3:b5):{3{a3}}))?((b1<=b0)>>(4'd2 * b1)):((b5?b0:a5)<{3{a2}}))}};
  assign y1 = ((6'd2 * (a0>p0))||((b5!=b0)|(-(-a4))));
  assign y2 = ((~&(a0<<<a4))&&(~&(-4'sd2)));
  assign y3 = $signed(($unsigned((p14?b1:b3))?(p7<<b3):{{p3,a2,b1}}));
  assign y4 = (!(((~^(a5|b1))-((a3<<<b4)<(-a5)))!=={(a1^~a4),(a0||a0),(b1==b2)}));
  assign y5 = ((+$unsigned(((|((a5?a1:a4)?$unsigned(a0):(~&a4)))^~(((a5/b1))^(^(~^b3)))))));
  assign y6 = {4{(2'd0)}};
  assign y7 = ((({3{p0}})-(5'd2 * p13))<{2{(p17&&p4)}});
  assign y8 = {3{((b5?a2:a4)===(b0?b0:b4))}};
  assign y9 = {2{(a2!==a5)}};
  assign y10 = (+(((a2)^~(-a5))?((a2?b5:b3)^(b3!=a5)):(~^(b5||b1))));
  assign y11 = (5'd5);
  assign y12 = {4{b3}};
  assign y13 = (|(^((-((b4>=a3)!=(a2<a1)))!==((b2-a3)^(~(-b4))))));
  assign y14 = ((b5<p5)<=(p15?b5:p8));
  assign y15 = {{(2'd1)},{(b1?p17:a0)}};
  assign y16 = (-a1);
  assign y17 = (-3'sd1);
endmodule
