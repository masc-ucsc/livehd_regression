module expression_00421(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(-2'sd1)}};
  localparam [4:0] p1 = (2'd3);
  localparam [5:0] p2 = ((5'd4)!=(3'd0));
  localparam signed [3:0] p3 = (((-3'sd2)?((5'sd11)?(5'd7):(2'sd0)):((3'd6)?(3'sd1):(-5'sd8)))?(((-4'sd7)?(-2'sd1):(-3'sd1))?(5'd17):(5'd28)):((5'd24)?(2'd0):(4'sd5)));
  localparam signed [4:0] p4 = (((2'd3)|(3'd1))!==((4'd15)^~(-3'sd3)));
  localparam signed [5:0] p5 = ((((4'sd3)<<<(4'd9))+((4'sd5)%(-4'sd1)))|(((4'd0)!=(-2'sd0))<<<((5'sd13)%(3'd5))));
  localparam [3:0] p6 = (4'd0);
  localparam [4:0] p7 = ((((-5'sd12)?(-2'sd0):(5'sd2))>>((4'sd5)?(3'd4):(3'd1)))>>>(|(~^({4{(3'd4)}}?((-2'sd1)>=(3'sd0)):((4'sd5)<(-4'sd2))))));
  localparam [5:0] p8 = ((((3'sd1)||(-3'sd2))<((4'd3)!=(2'd3)))=={4{(2'd3)}});
  localparam signed [3:0] p9 = {(2'd1),{1{{3{(-3'sd3)}}}}};
  localparam signed [4:0] p10 = ((!(2'd1))===(-5'sd6));
  localparam signed [5:0] p11 = ((^(&(^((3'sd0)<=(-4'sd0)))))<((^(5'd0))>=((3'sd3)<<<(5'd16))));
  localparam [3:0] p12 = (~(({(4'd2),(4'sd5),(-2'sd0)}<<{(5'd7),(4'd6),(4'd3)})?((6'd2 * (3'd4))?((-4'sd3)<(5'd8)):((5'd11)|(-4'sd7))):(+{1{(~&((4'd15)||(3'sd1)))}})));
  localparam [4:0] p13 = {{1{(3'sd3)}},((3'd7)>(5'd2)),((2'd3)+(4'sd2))};
  localparam [5:0] p14 = (-5'sd0);
  localparam signed [3:0] p15 = (~&(|((-3'sd0)||(4'sd6))));
  localparam signed [4:0] p16 = {4{((2'd0)<=(2'sd1))}};
  localparam signed [5:0] p17 = (~(5'd6));

  assign y0 = {a2,b4,a4};
  assign y1 = ({2{(a5|b4)}}&&((!(~^a4))>>$unsigned((a1-p5))));
  assign y2 = {2{{4{p16}}}};
  assign y3 = ({2{$unsigned(p16)}}?((p0&p8)>(p7<<p5)):((p5+a0)?(b0&&b1):{1{b3}}));
  assign y4 = (+{(^{(&(~|(~^(~|{a0,p5,p8})))),{{p14,p0},{{a4,p9,p13}}},{{p16,p1,p8},(~p6),(~&p11)}})});
  assign y5 = $unsigned((~&(+(p3?a1:p10))));
  assign y6 = (a2<<a3);
  assign y7 = ({1{(!{2{(p5!=p6)}})}}==((p8!=p12)|$signed((p7>p14))));
  assign y8 = ({{{p2,p17},(p4>=p7)}}&&{(p1&b3),{p10,p0},(p17==p11)});
  assign y9 = (({(+{a3})}===(5'd2 * (~a2)))&(~((p14<p12)^~(~&(!p11)))));
  assign y10 = ((3'd6)<<<(($unsigned(p14)=={1{a4}})));
  assign y11 = {1{b3}};
  assign y12 = ((b3<<<b3)+(a3==b3));
  assign y13 = ((a2>b4)*(b4===b4));
  assign y14 = ({p2,b1,a4}?{p4,p5,a5}:(p3<p9));
  assign y15 = ((~p13)&&(~p1));
  assign y16 = (5'd31);
  assign y17 = ((a1===b0)<<<(~^(a5>a2)));
endmodule
