module expression_00426(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{(-5'sd8)}}<(&((4'sd1)<=(3'd0))));
  localparam [4:0] p1 = (|{((5'd22)&&(-3'sd1)),((4'd3)!==(2'd0)),(-5'sd15)});
  localparam [5:0] p2 = {((-3'sd2)?(-5'sd12):(3'sd1)),{(5'd18),(2'd1)},(~|((-2'sd1)<(5'd29)))};
  localparam signed [3:0] p3 = {(((-2'sd1)?(4'sd0):(-5'sd0))?((3'sd1)?(2'd0):(-4'sd0)):{(5'd30)}),(((-5'sd1)?(2'd0):(4'sd5))?((3'd5)+(-4'sd3)):((2'd2)^~(3'd4))),({(4'sd0)}?((4'd11)>(5'd29)):((2'd2)<(3'd5)))};
  localparam signed [4:0] p4 = ((~^{{(-5'sd9),(3'd0),(5'sd1)},((4'sd7)?(4'd8):(-3'sd1))})>=({(5'sd13),(-3'sd2),(5'd11)}?(~&(4'd9)):(-5'sd10)));
  localparam signed [5:0] p5 = (3'd7);
  localparam [3:0] p6 = {2{(3'd4)}};
  localparam [4:0] p7 = {1{(-4'sd2)}};
  localparam [5:0] p8 = {({((3'd6)<<<(-4'sd1))}>>>((-5'sd15)<<(2'd0))),(!({(4'd5),(-2'sd0)}>>{(4'sd6),(3'd6)}))};
  localparam signed [3:0] p9 = {1{((-3'sd0)===(2'd3))}};
  localparam signed [4:0] p10 = (3'sd1);
  localparam signed [5:0] p11 = ({((5'd30)<(4'd13))}?{(-3'sd1),(4'sd4),(-5'sd11)}:((4'd8)?(3'sd3):(-4'sd7)));
  localparam [3:0] p12 = {4{(6'd2 * (2'd3))}};
  localparam [4:0] p13 = {((3'sd3)===(3'd3)),{(4'd2),(3'd0),(4'd4)},{((2'd0)<(4'd0))}};
  localparam [5:0] p14 = {1{((+((5'd26)?(2'd3):(5'sd10)))?((2'd2)?(3'd6):(4'd9)):((2'd1)?(-5'sd6):(4'd4)))}};
  localparam signed [3:0] p15 = (-(2'd3));
  localparam signed [4:0] p16 = ((((4'd8)^~(5'd6))|{4{(2'sd0)}})-({3{(4'd7)}}?(+(-4'sd2)):((5'd3)?(2'sd1):(2'd2))));
  localparam signed [5:0] p17 = (~&(!(2'sd1)));

  assign y0 = (-4'sd7);
  assign y1 = (((b0?a3:b0)<=(b5<b2))>((b2?b2:b4)?{4{a5}}:(b4!==b2)));
  assign y2 = $unsigned({1{((~|{2{p15}})&(~|(6'd2 * p0)))}});
  assign y3 = ((5'd2 * (3'd2))?{p1,p8,a5}:(b0?a0:p11));
  assign y4 = ((~^((p5==p8)+(p2&&p7)))^(-4'sd3));
  assign y5 = (~(-2'sd1));
  assign y6 = (~|(|(&(&{(~&$signed((-(4'd2 * {p14})))),(^((b0&b5)<={p17,p17,p11}))}))));
  assign y7 = {{3{$unsigned(p17)}},(3'd4),$signed($unsigned({{3{p5}}}))};
  assign y8 = ((a5%a2)/p8);
  assign y9 = (((a1==a5)>{4{p1}})?{3{(p9?p7:p9)}}:{((p9-p1)|(b0?p14:p17))});
  assign y10 = (-5'sd8);
  assign y11 = (&((p3>>p3)>(p16?p8:p17)));
  assign y12 = (~($signed($signed((|((-{p8,p13,p5})>>>((~^a1)>{a1})))))));
  assign y13 = ({a0,b0,p15}?(p6?b4:p7):(^b2));
  assign y14 = ((p12?b2:p4)?$signed((b4?b3:b0)):(a1?b2:p0));
  assign y15 = (~(+((!({a1,b3}|(&b0)))?{(a4?b0:a4),(p0>>p12),(~&a1)}:({a5,p11,b1}&{a1}))));
  assign y16 = $signed(((~^(-5'sd3))));
  assign y17 = (a5?p12:p1);
endmodule
