module expression_00061(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'sd0)&(3'sd0))&((5'sd0)&&(4'd10)))&&(~^((2'sd1)!==(4'sd1))));
  localparam [4:0] p1 = {3{{3{(2'sd1)}}}};
  localparam [5:0] p2 = (-{3{((&(4'sd3))^{4{(4'd6)}})}});
  localparam signed [3:0] p3 = {3{((5'sd14)&&(5'sd12))}};
  localparam signed [4:0] p4 = ((((2'sd0)<<<(2'd2))?(3'd5):(3'd7))?(((5'sd3)?(5'sd13):(-4'sd5))>>>(3'sd2)):((-5'sd3)&&((5'd5)*(2'sd0))));
  localparam signed [5:0] p5 = (|(4'd7));
  localparam [3:0] p6 = (-4'sd3);
  localparam [4:0] p7 = (({(5'sd4),(5'd3)}>{4{(3'd3)}})?(((4'd2)-(4'd5))>>>((5'sd5)==(4'd7))):(-5'sd8));
  localparam [5:0] p8 = (!(~(~(|((4'd14)!==(~^(4'd2)))))));
  localparam signed [3:0] p9 = (~|(((-2'sd0)?(4'sd2):(4'd1))?((3'sd1)&&(4'sd5)):((3'd7)?(-3'sd0):(-2'sd0))));
  localparam signed [4:0] p10 = (4'd11);
  localparam signed [5:0] p11 = {3{(((2'd1)>>(4'd5))>={1{(4'sd4)}})}};
  localparam [3:0] p12 = (~^((((-2'sd0)>(-3'sd3))?{(3'd1)}:((5'd31)<=(-5'sd2)))===(~|{(~|(2'd3)),((5'd23)?(3'sd3):(-2'sd0))})));
  localparam [4:0] p13 = {2{{4{(|(5'sd11))}}}};
  localparam [5:0] p14 = ({1{((^((2'sd1)-(5'd12)))^{3{(2'd2)}})}}!==({1{(&(4'd6))}}>=(-(!(5'd23)))));
  localparam signed [3:0] p15 = (4'd2 * ((2'd2)!==(3'd3)));
  localparam signed [4:0] p16 = {4{{4{(5'd25)}}}};
  localparam signed [5:0] p17 = {{{{(5'd24),(3'd4)},((5'd3)|(5'd14)),(6'd2 * (2'd0))},{{3{(2'd3)}}},({(5'sd3)}<<<((3'sd0)|(-2'sd1)))}};

  assign y0 = (($signed(a2)^(p5<<b3))^~{{b1},(a2?p9:a4),(a0^p17)});
  assign y1 = (-3'sd3);
  assign y2 = {2{$unsigned(((b3===b5)^(a3)))}};
  assign y3 = (((a5*a4)>>(b0||a3))>>((b4!=b2)<(a5!==a3)));
  assign y4 = ((3'sd3)^((2'd1)<<<{(~&p8),(4'd2),{p0}}));
  assign y5 = (3'd2);
  assign y6 = ({((4'd1)+(3'sd3)),((a2?b0:b4)!=(b2)),(2'd3)});
  assign y7 = (-2'sd1);
  assign y8 = {{(p4?a5:p8),(a3?a4:b2)},({a2,b4,a2}?(b4?a3:b5):(p13?a3:a5))};
  assign y9 = (((3'd6)&(~a1))-(4'd6));
  assign y10 = (2'd0);
  assign y11 = (2'd2);
  assign y12 = $unsigned((-5'sd8));
  assign y13 = {2{(6'd2 * {2{p6}})}};
  assign y14 = {((2'd1)&&((b2?a2:a1)?(&(!b3)):(a2?a1:a3)))};
  assign y15 = (({4{b4}}^(p10?b4:b4))<$unsigned((4'd2 * $unsigned(a5))));
  assign y16 = {{(!(p12)),(b5===a3),(p8<p11)},(((a4^b1)<<<(b1!==b5))>>>{2{{4{p14}}}})};
  assign y17 = ((-b1)<<<(4'd10));
endmodule
