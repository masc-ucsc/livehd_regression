module expression_00448(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(+(~^{(5'd26),(-5'sd9)})),{{2{(5'd21)}}}};
  localparam [4:0] p1 = (~&((~|(4'd3))^((-3'sd2)?(5'd9):(4'd5))));
  localparam [5:0] p2 = ({{(4'd2),(5'd26)}}|(|(~&{(4'sd4),(-4'sd4)})));
  localparam signed [3:0] p3 = (2'sd1);
  localparam signed [4:0] p4 = (((5'sd6)?(5'd21):(4'sd2))?(5'd2 * {3{(3'd5)}}):((4'd3)?(-5'sd12):(3'd4)));
  localparam signed [5:0] p5 = ((((5'sd11)?(4'd9):(2'd3))?(~&(4'sd2)):(-(-4'sd7)))?((+(5'd12))?((-5'sd11)>>(3'd7)):{(5'd12)}):(((-2'sd0)<<<(3'sd3))^~{(5'd6),(4'd13),(3'sd2)}));
  localparam [3:0] p6 = {2{(((-3'sd2)^~(5'd9))^~(-(3'd2)))}};
  localparam [4:0] p7 = (+(!(((2'd0)>=(5'd1))<(~&(4'sd5)))));
  localparam [5:0] p8 = (-{({{(-2'sd1),(5'sd9)}}=={(-3'sd0),(2'd3),(5'd8)}),{3{(~|(4'd10))}}});
  localparam signed [3:0] p9 = {(((2'sd0)|(-3'sd2))<<(~|((-4'sd5)&&(4'd2)))),(((5'd22)>>(5'sd8))<<<((2'sd0)?(-3'sd1):(5'sd6)))};
  localparam signed [4:0] p10 = {({(-3'sd1),(2'd2),(4'sd1)}+((4'd14)?(-3'sd3):(-4'sd4)))};
  localparam signed [5:0] p11 = {3{{1{(~|(5'sd2))}}}};
  localparam [3:0] p12 = {((3'd2)>>>(5'sd8))};
  localparam [4:0] p13 = (^(!((-5'sd15)>(2'sd1))));
  localparam [5:0] p14 = ((4'sd7)?(2'd2):(4'd0));
  localparam signed [3:0] p15 = (5'd22);
  localparam signed [4:0] p16 = {{(2'sd1),(4'd2),(3'd0)}};
  localparam signed [5:0] p17 = (5'd29);

  assign y0 = (((a1<a5)>>>(p5<<<p11))||(4'd2 * (p2?a0:p14)));
  assign y1 = (((4'sd2)&&(b0<<a3))!==((a5^~b2)<<{b1,b2,b4}));
  assign y2 = $unsigned($signed(((a2?a2:b0)?(~|b4):(3'd7))));
  assign y3 = ((b2?p15:b0)^((5'd2 * a0)^(b1&&b5)));
  assign y4 = {4{a3}};
  assign y5 = {(p16^~b5),{1{(3'd4)}}};
  assign y6 = (-(3'sd3));
  assign y7 = {4{(({b0}))}};
  assign y8 = (((b3?p8:p9)?(p11<b5):(a2!==b3))|((p16?b1:b0)/p7));
  assign y9 = {2{p9}};
  assign y10 = $unsigned((($signed(p13)?{p4}:{p15})));
  assign y11 = (2'd3);
  assign y12 = ((~&(b1>>b5))^((p0-p5)&(~^p4)));
  assign y13 = {{(p16?p11:b0),(p11?p11:p17)},(({p15}?$signed(p10):(!p5)))};
  assign y14 = (-b3);
  assign y15 = ((2'd2));
  assign y16 = ($signed($unsigned((|(+(2'd1)))))^~(4'd7));
  assign y17 = (5'd28);
endmodule
