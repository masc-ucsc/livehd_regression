module expression_00907(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{2{{2{{3{(4'd15)}}}}}}}};
  localparam [4:0] p1 = (~|((4'sd0)||(2'sd0)));
  localparam [5:0] p2 = {2{((-2'sd0)?(-4'sd4):(4'sd2))}};
  localparam signed [3:0] p3 = (4'd9);
  localparam signed [4:0] p4 = ((2'd2)^((3'sd3)>>>(4'd4)));
  localparam signed [5:0] p5 = ((((2'd1)?(5'd12):(3'd6))|{(-5'sd9)})?(^{1{((-5'sd5)?(5'sd3):(3'd7))}}):({(5'd27),(2'd3),(3'd3)}<<(4'd2 * (5'd19))));
  localparam [3:0] p6 = (((4'd7)?(5'd23):(2'd0))?{1{(+(2'd3))}}:((4'sd4)?(3'sd0):(2'd1)));
  localparam [4:0] p7 = ({{(-3'sd2),(2'd0),(-4'sd0)},(~{1{(4'sd5)}})}<<<(^(~^(+((2'd2)>>(4'd4))))));
  localparam [5:0] p8 = {4{((2'd2)>>(2'd1))}};
  localparam signed [3:0] p9 = (~^(^(-{4{((5'sd9)?(5'd21):(2'd3))}})));
  localparam signed [4:0] p10 = (-5'sd12);
  localparam signed [5:0] p11 = ({4{(2'd1)}}+(^((3'sd0)<(-4'sd0))));
  localparam [3:0] p12 = {3{((2'd2)==(3'sd2))}};
  localparam [4:0] p13 = (((|(-5'sd10))>=(|(4'd10)))<(~((-2'sd1)/(2'sd1))));
  localparam [5:0] p14 = (&(~&((!(5'd27))?((5'd2)?(-3'sd0):(2'd1)):((4'd13)?(2'd2):(-2'sd0)))));
  localparam signed [3:0] p15 = (((-3'sd1)?(-4'sd3):(2'd1))?((5'd2)+(5'sd2)):((4'd1)?(3'sd2):(3'sd3)));
  localparam signed [4:0] p16 = ((((3'd0)+(-2'sd0))===((4'd6)^(5'sd6)))?{(~^((5'd18)?(2'd2):(3'sd1)))}:{(((3'd5)?(4'sd3):(4'd0))^(&(5'd18)))});
  localparam signed [5:0] p17 = {(5'sd7),(5'd15),{{3{(-2'sd1)}}}};

  assign y0 = ((((a1&a5)^~(b4==b3))!==((5'd2 * b1)&&(a3===b2)))===((a2-b5)*(b1!==b4)));
  assign y1 = (~&(~(!(&(!b1)))));
  assign y2 = (-2'sd0);
  assign y3 = (~^{3{p0}});
  assign y4 = $unsigned({(&(|p3)),(~^(~a1))});
  assign y5 = {3{(^a1)}};
  assign y6 = ((~&(~{a4,p14,p13}))?((5'sd8)?(5'd7):(2'sd1)):(~((b2?p11:p6)<(2'd0))));
  assign y7 = {3{(2'sd0)}};
  assign y8 = {4{(p16&b0)}};
  assign y9 = ((a0?a5:a3)^(+(b5>a5)));
  assign y10 = (((a1?p17:p14)?{4{p5}}:(4'd10))<<<{1{((3'd7)|(-p10))}});
  assign y11 = ((-((-3'sd1)?(p10?p6:p2):(5'd19)))<=(+(4'd1)));
  assign y12 = ((a2|a4)<(b5?b5:a1));
  assign y13 = ((5'sd2)>=((p9>>a0)|(a3-p1)));
  assign y14 = ({1{$unsigned(p10)}}>=(-2'sd0));
  assign y15 = {{(p3<p13),(a1?a0:a4)},((b0?p2:p15)&(4'sd2)),({(3'd5)}>>>(-4'sd2))};
  assign y16 = (4'd2 * (3'd6));
  assign y17 = (^(+((a0>a1)>=(a5?b4:b5))));
endmodule
