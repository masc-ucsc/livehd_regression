module expression_00320(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{2{(3'd3)}},(&{1{(-5'sd2)}})};
  localparam [4:0] p1 = ({3{(-4'sd6)}}?((5'd16)?(2'd0):(2'd2)):((2'd1)?(4'd1):(-5'sd10)));
  localparam [5:0] p2 = (((-2'sd0)&&(-4'sd0))^((5'd0)&(4'd13)));
  localparam signed [3:0] p3 = (5'd25);
  localparam signed [4:0] p4 = (!{1{(~^((3'd6)!=((2'd1)==(5'd21))))}});
  localparam signed [5:0] p5 = (((3'd4)?(2'sd1):(4'sd5))?{(5'sd9),(3'd3),(3'd5)}:(~&(3'sd2)));
  localparam [3:0] p6 = ((3'd4)||(3'd3));
  localparam [4:0] p7 = (-2'sd0);
  localparam [5:0] p8 = ((4'sd0)&&(|(5'd27)));
  localparam signed [3:0] p9 = (3'd5);
  localparam signed [4:0] p10 = ({4{(-3'sd1)}}>>>({4{(-5'sd2)}}!={4{(5'sd6)}}));
  localparam signed [5:0] p11 = {2{{(3'd2),(-5'sd2),(5'd30)}}};
  localparam [3:0] p12 = ((((2'sd0)==(-2'sd1))?((-3'sd3)?(5'd25):(4'sd1)):{(3'd3),(2'd1)})<<{{{(2'd2),(2'd3)},((-3'sd0)||(2'sd0))}});
  localparam [4:0] p13 = (~|(2'd0));
  localparam [5:0] p14 = {2{{3{(5'd14)}}}};
  localparam signed [3:0] p15 = (((-2'sd1)<((-3'sd2)+(2'd1)))>>>{1{(3'sd3)}});
  localparam signed [4:0] p16 = (({4{(-5'sd10)}}^~(-3'sd3))^((6'd2 * (3'd3))+(-2'sd0)));
  localparam signed [5:0] p17 = {((2'sd1)?(3'sd3):(5'd16)),{((5'd26)&(2'sd0))},(-5'sd10)};

  assign y0 = ({1{(({1{{4{a0}}}}-(2'sd1)))}});
  assign y1 = {2{(p2?p8:p13)}};
  assign y2 = {(-{{({(-b4)}||(-(-p12))),{{(!(p2||p11))}}}})};
  assign y3 = (((~&(p6<<p4))>>>(p8!=a5))>>((b4!=a2)!=(p14|p9)));
  assign y4 = (5'd2 * b2);
  assign y5 = (-4'sd2);
  assign y6 = (((p8>b4)&&(p14?p12:b2))?{3{a0}}:(~^(~|(&b4))));
  assign y7 = (((4'd2 * (a0&a0)))<=(~&(+$signed($signed((a3+b0))))));
  assign y8 = $signed(($signed(b4)^(a3)));
  assign y9 = ({p17}?{a1}:(b1?a3:p10));
  assign y10 = $unsigned((p5?p9:p10));
  assign y11 = {{{p6,p15},(a1!==a2)},({a5,a4,a4}!==(a1!=a1))};
  assign y12 = {3{(p16?p15:a1)}};
  assign y13 = ((((5'sd2)===(b5<<b4)))||(|$unsigned(((-3'sd1)<<<{p15}))));
  assign y14 = {{{p4,p6}},{(p13&p8)}};
  assign y15 = {(a5?a3:p14),(~^(p9?b3:a0)),({1{p5}}^{1{a0}})};
  assign y16 = (~^((((~a1)!=(a4<<<a2))<=((p3^~p8)))||$unsigned($unsigned(((a3^~p16)&(p0<=p8))))));
  assign y17 = $unsigned(p4);
endmodule
