module expression_00128(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{((3'd5)|(5'd8))}}>>>(2'sd1));
  localparam [4:0] p1 = ((3'sd2)!=(2'd2));
  localparam [5:0] p2 = ((-4'sd5)?(2'd2):(-4'sd7));
  localparam signed [3:0] p3 = (({(5'd2 * (2'd3))}^~((5'sd4)<<<(2'sd1)))<=({(-3'sd3),(4'd7),(3'd7)}<<{{(2'd0),(-2'sd1)}}));
  localparam signed [4:0] p4 = ({(3'd3),(4'd10),(-3'sd0)}!==(~&(4'd4)));
  localparam signed [5:0] p5 = ((6'd2 * (6'd2 * (5'd30)))||(((3'd1)-(5'sd0))==(-3'sd2)));
  localparam [3:0] p6 = (~^{((!(2'd1))&(~|(5'sd6))),(((3'd7)||(5'd7))<<<{(2'sd0),(3'd7),(3'd0)})});
  localparam [4:0] p7 = {((2'sd1)>((2'sd0)>>(4'd5))),{(~{(2'sd0)}),{(4'd2),(4'd0)}}};
  localparam [5:0] p8 = {2{(~^(2'd0))}};
  localparam signed [3:0] p9 = (^(+(((5'sd1)==(~(4'sd0)))-(|{1{{1{(~|{3{(3'sd0)}})}}}}))));
  localparam signed [4:0] p10 = ({3{(3'd6)}}^{3{(4'd0)}});
  localparam signed [5:0] p11 = {({((-2'sd0)!=(-5'sd7)),{((5'd31)?(-2'sd0):(-4'sd3))}}==({(4'd13),(5'sd9),(5'd12)}?((2'd2)?(4'd6):(5'd8)):{(5'd9)}))};
  localparam [3:0] p12 = (~&(!(^({{2{{(2'd2),(2'd1),(2'd0)}}}}^{3{(^(5'd29))}}))));
  localparam [4:0] p13 = (~{(3'd6),(-2'sd0)});
  localparam [5:0] p14 = (&((3'sd2)==(4'sd1)));
  localparam signed [3:0] p15 = (((~|(2'sd1))===((-4'sd0)^~(-5'sd6)))===(((5'd4)^~(3'sd2))&((5'sd2)>(3'd4))));
  localparam signed [4:0] p16 = (~(+(~^(2'd0))));
  localparam signed [5:0] p17 = {3{((-3'sd2)+(4'sd6))}};

  assign y0 = (~&{3{(!p1)}});
  assign y1 = {4{$signed((p2^a3))}};
  assign y2 = {(+(5'd9))};
  assign y3 = (5'd2 * (2'd3));
  assign y4 = {((a5?a1:p14))};
  assign y5 = (~|(&(!((+(|({3{p8}}?{4{p12}}:(-p17))))>>((p14?b0:p9)<=(p9?p12:p4))))));
  assign y6 = (4'sd4);
  assign y7 = (^{(2'd0)});
  assign y8 = ((((p2==a0)!=(b1<<p4))^((b4<b3)!==(a5>=a0)))>(((p8/p13)>(b1===a1))^((p11>>a1)&&(b5>=p13))));
  assign y9 = (-p13);
  assign y10 = (4'd2 * {{p6,p12,p0}});
  assign y11 = {2{$unsigned((~|((~a4)==(+a5))))}};
  assign y12 = (((a2>>>p9)?(b3?a2:b5):(b0?a1:b0))?{2{{1{(b3?a2:p5)}}}}:((a0?p0:p11)||(p1>=p2)));
  assign y13 = (({4{p10}})<=(5'sd15));
  assign y14 = $signed(p7);
  assign y15 = ((&((b0<<b0)?(b3<<<p10):{1{b3}}))?(~((5'sd3)===(3'd1))):((4'sd3)==(p3<<<b2)));
  assign y16 = (~^(~|(((p1^p17)==(p17+p15))?(p2?a1:p13):{(b0>a0),(~&p1)})));
  assign y17 = ((|(4'd2 * a1))?(~(2'd3)):(p15?p14:b3));
endmodule
