module expression_00897(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(((~(4'd3))<<(-(-5'sd7)))<=(((-4'sd3)<=(5'd25))<(~(2'sd0)))));
  localparam [4:0] p1 = (4'd7);
  localparam [5:0] p2 = (~|{(~|((-4'sd5)?(5'd12):(-4'sd7))),(-(4'd10))});
  localparam signed [3:0] p3 = (-2'sd0);
  localparam signed [4:0] p4 = ((2'd1)?(5'd24):(5'd11));
  localparam signed [5:0] p5 = ((-{(&(5'd14)),(~|(2'd1)),{(4'd8),(-5'sd5)}})+({(-3'sd0),(-2'sd0),(4'd10)}>{4{(5'sd8)}}));
  localparam [3:0] p6 = {2{(((2'd1)===(4'd1))!=(&{3{(4'd11)}}))}};
  localparam [4:0] p7 = (~&(+(((5'd29)?(-3'sd2):(-2'sd1))>>(+(3'sd2)))));
  localparam [5:0] p8 = ((~&({(3'd4),(3'd4),(-5'sd12)}>>>(|(5'd14))))<(3'd2));
  localparam signed [3:0] p9 = (^((3'd1)|(5'd21)));
  localparam signed [4:0] p10 = (!(~((2'd2)^(!((~(2'sd1))?((4'd8)?(2'd2):(2'd3)):(|(2'sd0)))))));
  localparam signed [5:0] p11 = {2{(~&(^(4'd7)))}};
  localparam [3:0] p12 = (((5'd27)<=(-4'sd2))&((5'd0)>>(5'sd10)));
  localparam [4:0] p13 = {((2'd2)?(3'sd1):(3'sd1)),(((3'sd2)?(2'd0):(3'sd0))>>>((3'sd0)<<<(3'd2)))};
  localparam [5:0] p14 = (-2'sd1);
  localparam signed [3:0] p15 = ((+(3'd5))?{2{(4'd1)}}:{3{(2'sd1)}});
  localparam signed [4:0] p16 = (^(5'sd3));
  localparam signed [5:0] p17 = (^(~&(~&(((~&(2'd3))!=((4'sd3)*(-3'sd1)))&(-((4'd11)<<<(5'd17)))))));

  assign y0 = (((p5%p14)>=$signed(p5))?(4'd2 * (p2?p2:p13)):(p12?p5:p8));
  assign y1 = (a5-p9);
  assign y2 = (-5'sd3);
  assign y3 = ($signed(((a0<a0)>>(b1>>>a5)))+($unsigned((!(^b4)))<<((b0*a4)>>>(~^b3))));
  assign y4 = ($signed(a1)===$signed(b3));
  assign y5 = ((!{(a0?a0:b2)})^((~a3)^(b2?b2:p13)));
  assign y6 = (3'sd0);
  assign y7 = (((b5+b0)===(b2|b5))&&({(a1||a5)}!==(a5>>b5)));
  assign y8 = (4'sd2);
  assign y9 = ((!(~^((4'd12)!=(3'd5))))<(-2'sd0));
  assign y10 = ((&{({p2,p15,p3}?{p0,a5}:(+b2))})<((~&{p8,p0})?(b1&p10):(p17<=b2)));
  assign y11 = (~({(~&{((~|a3)),(-(b4<=a3))})}!==((a1&&a2)?(b5>=b3):$unsigned({2{a4}}))));
  assign y12 = (3'sd1);
  assign y13 = {{b1,a2},(3'd4),$unsigned($signed(b3))};
  assign y14 = ((((((p16?p6:p14))=={p11,p7,p3})))>>>(({p17,p2}>(p7?p0:p0))!={(p2?p7:p11)}));
  assign y15 = ({((p13||p6)?(b2>>a1):(p17?a5:a2))}>>>{(b3>=a3),(a5!==a0),(b0?a0:b2)});
  assign y16 = (|(((p3^~p13)>=(p4==a1))|((p1>>a0)==(~|(p4%p8)))));
  assign y17 = ((p0<<p1)%p10);
endmodule
