module expression_00569(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(|((-(3'd0))!==((4'sd6)!=(5'sd3))))}};
  localparam [4:0] p1 = (((5'd20)?(5'd19):(4'd10))<(|((-4'sd3)&(5'd29))));
  localparam [5:0] p2 = ((-3'sd2)^~(2'sd1));
  localparam signed [3:0] p3 = {{1{{2{(((5'sd5)||(-3'sd2))<<{3{(2'd3)}})}}}}};
  localparam signed [4:0] p4 = (+(~|((^(5'd0))?((4'd13)?(-5'sd9):(2'd1)):(4'd1))));
  localparam signed [5:0] p5 = ((((6'd2 * (2'd0))>>>((2'd1)?(-3'sd3):(-5'sd8)))>(~(-((-2'sd1)?(-3'sd1):(-2'sd0)))))>((!(-3'sd2))?(3'd0):(~|(3'sd1))));
  localparam [3:0] p6 = (~^{(({(2'd3)}<{(-3'sd0),(3'd5),(-5'sd7)})<<({(-4'sd7)}&((4'd4)?(5'sd13):(-2'sd0))))});
  localparam [4:0] p7 = (~^(-4'sd3));
  localparam [5:0] p8 = (((4'd12)?(5'd10):(5'd0))?(~(4'sd4)):((4'sd5)?(-2'sd0):(-4'sd0)));
  localparam signed [3:0] p9 = {({3{(-5'sd5)}}<<((5'd22)?(5'sd4):(4'd12))),(((2'sd0)?(3'sd0):(-4'sd6))?((-3'sd1)?(2'd1):(5'd28)):{(5'd17),(4'd13),(3'd7)})};
  localparam signed [4:0] p10 = {{(2'd1),(3'd2),(3'd3)},{4{(-2'sd0)}},{(-3'sd1),(3'sd0),(3'sd3)}};
  localparam signed [5:0] p11 = ((2'sd1)<=(((2'd2)>=(5'sd4))?((3'd7)>=(5'd8)):((2'd3)>>>(-2'sd0))));
  localparam [3:0] p12 = ((((3'd4)<=(4'sd0))&&(2'd1))-{2{((2'sd1)^~(3'd2))}});
  localparam [4:0] p13 = {2{(5'sd12)}};
  localparam [5:0] p14 = {1{(((5'd2)>=(5'd7))!==((-3'sd3)!=(4'd6)))}};
  localparam signed [3:0] p15 = (5'sd10);
  localparam signed [4:0] p16 = (~|(~{1{(^(-4'sd3))}}));
  localparam signed [5:0] p17 = (({1{(-5'sd6)}}==((2'd2)<<(2'd2)))|{2{((5'd2)!==(4'd7))}});

  assign y0 = (((b1&p4)&{3{p3}})?{3{(6'd2 * b1)}}:{2{(p12==p0)}});
  assign y1 = (!(($unsigned((p11!=b5)))-(~|((5'd11)&(-2'sd1)))));
  assign y2 = (&(-4'sd6));
  assign y3 = ((~|(p6))?{p1,p15,p5}:(+{a3}));
  assign y4 = ({4{p8}}&(b4!==b1));
  assign y5 = ({2{((+p10)|{4{p17}})}}>>>(|({1{(p2>>p4)}}-(p13>p0))));
  assign y6 = {3{{4{p16}}}};
  assign y7 = (^($signed(((p13+p15)>>(p9*p0)))^~$unsigned((((p14==a1)&(a4|p10))))));
  assign y8 = (5'd15);
  assign y9 = (2'd2);
  assign y10 = ((~&(p16==p1))?((p12)<=(p9?p0:p17)):($unsigned(p10)|(5'd16)));
  assign y11 = $unsigned((4'd4));
  assign y12 = (!(~(-2'sd0)));
  assign y13 = (a3?b0:p15);
  assign y14 = (p3?p11:p4);
  assign y15 = (4'd14);
  assign y16 = ((b2<p2)?$signed(b0):(p8?p0:p11));
  assign y17 = (&(3'sd1));
endmodule
