module expression_00467(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd30);
  localparam [4:0] p1 = ({3{(3'd2)}}?((5'sd10)>(-3'sd2)):((4'sd7)+(2'd3)));
  localparam [5:0] p2 = ((3'sd3)?(((3'sd1)?(3'sd0):(4'd15))^~(4'd14)):(^(|(~(-4'sd7)))));
  localparam signed [3:0] p3 = ((((-5'sd5)^(4'd10))==(5'sd4))!==((3'sd0)?(-3'sd0):(2'd1)));
  localparam signed [4:0] p4 = ((-2'sd1)|(-2'sd0));
  localparam signed [5:0] p5 = (+(|((-(3'd1))+((4'd2)^~(3'd7)))));
  localparam [3:0] p6 = (((-3'sd0)>=(-5'sd1))>((3'sd3)/(-2'sd0)));
  localparam [4:0] p7 = (~(!(((2'd0)>=(-5'sd9))>=((5'sd8)^~(5'd10)))));
  localparam [5:0] p8 = ({2{(|(~&(3'd1)))}}<<<(~(&((|(5'd16))>>>{3{(-3'sd1)}}))));
  localparam signed [3:0] p9 = (6'd2 * (~(3'd4)));
  localparam signed [4:0] p10 = ({(((4'd3)>>(3'sd1))!=((5'd3)>(4'sd1)))}<({{(-4'sd5),(4'd0),(-5'sd0)},(3'd5)}>>>(3'd5)));
  localparam signed [5:0] p11 = {3{((!(4'd10))&&((3'sd2)!==(-4'sd2)))}};
  localparam [3:0] p12 = {2{((3'd6)+(-4'sd5))}};
  localparam [4:0] p13 = ((4'd5)?(5'sd13):((3'd5)|(2'sd1)));
  localparam [5:0] p14 = ({{(-4'sd4),(4'sd7),(5'sd0)},((-3'sd1)?(-4'sd2):(4'd8))}^~(((3'd4)?(-5'sd8):(5'd20))+((-4'sd0)?(-4'sd5):(5'd24))));
  localparam signed [3:0] p15 = ((-5'sd4)&(((-3'sd2)!==(-5'sd12))<=(!(5'd25))));
  localparam signed [4:0] p16 = (-{2{{4{(5'd9)}}}});
  localparam signed [5:0] p17 = ((((3'sd3)==(5'd30))<=((5'd20)?(5'sd2):(3'd4)))<=(((4'd15)<<(3'sd2))?((4'sd5)<<(2'd0)):((2'd1)>=(4'd6))));

  assign y0 = ((&(~^p15))?(~^(p10+a3)):{(p13?p8:p14)});
  assign y1 = $unsigned(((a3?a4:a0)>=((b3==p4)^$signed(p6))));
  assign y2 = ((((~&a1)==(&b3))==(~&(&(a2^~b3))))!=(((~|p17)<(!p10))>>((b1&b4)?(b4|b4):(&p1))));
  assign y3 = $signed($unsigned({((b5^a2)?(b5>=a2):{p7,a1,p2}),((a1?b1:p2)?$signed(p2):$signed(p12)),((p3!=p5)?$signed(p8):(6'd2 * p2))}));
  assign y4 = (4'sd4);
  assign y5 = ((~^(+(~^b1)))?{1{(-(~b0))}}:{1{(a0?p2:a4)}});
  assign y6 = ((-3'sd3)^(~|a4));
  assign y7 = (~&$unsigned(({2{$signed((a3?a0:b4))}}===(~((a5>a4)>>(b3?b2:b1))))));
  assign y8 = (3'd1);
  assign y9 = ((a5!=a4)&&(b0?a3:b0));
  assign y10 = (|{2{(~|(((&p8)|(p14^a3))&((b4|p3)==(a4!=p3))))}});
  assign y11 = (b3?b4:a0);
  assign y12 = $unsigned(b1);
  assign y13 = ($signed(((~(p3-p9))==(p9&b1)))==(&($unsigned(p15)?(a1?p5:p5):$unsigned(p2))));
  assign y14 = (^{1{b4}});
  assign y15 = (p12?b2:p6);
  assign y16 = (((!{4{a2}})>>>(p3?p7:b0))||((b5+a0)>=(b1>=a0)));
  assign y17 = ((((4'd2 * a1)<<(b4?a1:a1))!==(a5?b5:a3))>((a1?a1:a4)==((~^b1)^~(b0|p0))));
endmodule
