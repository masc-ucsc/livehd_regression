module expression_00602(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({((5'd28)?(2'd2):(2'sd0)),((-2'sd1)?(2'd3):(3'd1))}?((4'sd0)?(-5'sd13):(-3'sd3)):(((-5'sd6)?(3'd3):(4'd7))==(-(2'd0))));
  localparam [4:0] p1 = (-{(-2'sd0)});
  localparam [5:0] p2 = {(!((2'd3)?(5'd27):(-5'sd15))),{(2'd0),(3'sd1),(4'd3)}};
  localparam signed [3:0] p3 = ((4'd2)===(5'sd9));
  localparam signed [4:0] p4 = (!{4{(5'd30)}});
  localparam signed [5:0] p5 = (({(5'sd8),(4'd7)}&&(~|(4'd13)))?{2{(^(4'd10))}}:{3{((3'sd1)||(5'sd1))}});
  localparam [3:0] p6 = ((2'd2)?((-2'sd0)*(5'd2)):((2'd2)/(2'sd1)));
  localparam [4:0] p7 = ((3'sd2)|{{{(4'd13),(5'd24)},(3'd3),(5'd4)}});
  localparam [5:0] p8 = (4'd1);
  localparam signed [3:0] p9 = (-(5'sd9));
  localparam signed [4:0] p10 = (|((2'd1)?(4'sd6):(2'd0)));
  localparam signed [5:0] p11 = {1{({4{(2'sd0)}}<(((5'sd15)<=(4'd9))>>{2{(5'sd3)}}))}};
  localparam [3:0] p12 = {3{({3{(5'd9)}}<=((5'd18)<<(3'sd2)))}};
  localparam [4:0] p13 = ((4'd3)!=(4'd11));
  localparam [5:0] p14 = ({2{(^(3'sd2))}}!={3{((-2'sd0)!==(-5'sd11))}});
  localparam signed [3:0] p15 = (!{(-(2'sd1))});
  localparam signed [4:0] p16 = (-3'sd0);
  localparam signed [5:0] p17 = (3'sd0);

  assign y0 = {3{{4{a4}}}};
  assign y1 = (~|$unsigned((4'd10)));
  assign y2 = (((((b1<=a0)>(a3^~b1))!==$unsigned((5'd2 * a1))))<=($unsigned(((-5'sd3)))));
  assign y3 = (5'd2);
  assign y4 = (!(|(+(!(-((!(|b4))/b0))))));
  assign y5 = {(p13>>p11),(~(b1>>>p2))};
  assign y6 = ((p11||a4)||(2'sd0));
  assign y7 = {4{{1{{p0,p8,p17}}}}};
  assign y8 = {2{{3{(a2?b5:b5)}}}};
  assign y9 = ((p4|p7)>(a1&&p3));
  assign y10 = (&$unsigned((((a2/b1)?(a0?a5:a0):(p4?p8:p7))-((~|((b4)))==((a1>>>p9)>>>(p11*b0))))));
  assign y11 = (5'd16);
  assign y12 = ({1{({4{p12}}+(3'd2))}}<(4'd15));
  assign y13 = (a3!==a2);
  assign y14 = $unsigned((({4{b4}}==((&a3)>(a1?a0:a4)))!==((~^(-(b3)))|($unsigned(a1)>(b0^a3)))));
  assign y15 = ({(p1&&b3),{a3,a0}}<=({b5,a4,b3}-(a3&&p11)));
  assign y16 = $unsigned({$unsigned((5'sd6)),((b5?b1:p9)?(p8?p5:a4):(p3?p2:b4))});
  assign y17 = (b4?p5:b0);
endmodule
