module expression_00778(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(~((&((-2'sd0)==(5'd3)))-(+((2'd1)<=(5'd18))))));
  localparam [4:0] p1 = (^(^({(5'd9)}+{(4'd7),(4'd5)})));
  localparam [5:0] p2 = ((((2'd3)?(2'd3):(2'd2))?{(3'd0),(2'd1)}:((3'd4)?(2'sd1):(2'd3)))?({(5'sd5),(2'sd0),(-2'sd1)}>>>((-2'sd1)|(5'd7))):(((5'sd11)&&(-4'sd3))?{(-4'sd5)}:((-3'sd2)>>(5'd7))));
  localparam signed [3:0] p3 = ({2{(5'sd10)}}?((-2'sd1)!==(5'sd1)):((3'd0)>>(3'd1)));
  localparam signed [4:0] p4 = (4'd10);
  localparam signed [5:0] p5 = {((+(4'sd1))||((2'd3)>=(2'd2)))};
  localparam [3:0] p6 = {{1{(-4'sd4)}},(~|(5'd1)),(&(2'd2))};
  localparam [4:0] p7 = (^(!{1{{2{(5'd0)}}}}));
  localparam [5:0] p8 = {((~(((3'd7)^~(-2'sd0))?((-2'sd0)&&(3'sd2)):((-4'sd1)-(-4'sd5))))-(~&({(4'd15),(2'd2),(2'd2)}?{(-2'sd0),(-3'sd3)}:((3'd4)?(-5'sd8):(2'sd1)))))};
  localparam signed [3:0] p9 = (!(4'd1));
  localparam signed [4:0] p10 = (&(!((2'sd1)?(4'sd0):(4'd8))));
  localparam signed [5:0] p11 = ((!(-4'sd7))<<(2'd0));
  localparam [3:0] p12 = (((2'd3)?(2'd2):(5'sd13))?(~&((3'd1)&&(4'd0))):(-(!((-3'sd3)?(4'd12):(2'd1)))));
  localparam [4:0] p13 = {{2{(4'd14)}},{2{(3'sd0)}}};
  localparam [5:0] p14 = (!(~^{3{(~(5'd31))}}));
  localparam signed [3:0] p15 = {3{(5'd2)}};
  localparam signed [4:0] p16 = (5'd30);
  localparam signed [5:0] p17 = ((-5'sd6)?(2'd0):(5'd20));

  assign y0 = {(p10==p10),{p11,p16,p1},{(!p6)}};
  assign y1 = (a4!==a0);
  assign y2 = ((~|{$signed((p12^a1))})^~(&$signed((b4?b1:p6))));
  assign y3 = (b4&b5);
  assign y4 = ({4{(a1<p3)}}?((|(p16?b0:p1))<<<{1{(p2?p9:a5)}}):(!(^{4{p7}})));
  assign y5 = (((b4<a5)>>(a3&b5))!==(~&((b2|a1)!==(a2==a3))));
  assign y6 = ({1{{2{((a3==b2)===(b0!=b3))}}}}^({4{p4}}<<<({1{a3}}<<<(a3!==b1))));
  assign y7 = (~|(-((|((a5<<b4)>=(~|a4))))));
  assign y8 = (((~&(~^p14))==(|(p4|p10)))>>(~|(&(6'd2 * (~&(~&p14))))));
  assign y9 = (~^((p7?p7:b3)?(+($unsigned(b1))):$signed((!{b5}))));
  assign y10 = (((~&b5)?(~b5):(|p8))?(+(~|(^(b0?p1:b5)))):((-p17)?(^b3):(b0?b5:a4)));
  assign y11 = (+(~|(((p1-p7)!=(p6>>b1)))));
  assign y12 = (~&({1{a2}}==(~&a4)));
  assign y13 = (5'd4);
  assign y14 = (&p17);
  assign y15 = (((b1^~b5)?(-b0):(a5?b4:b4))||{(5'd31),(a0+a0),(a3&a5)});
  assign y16 = $signed({4{b5}});
  assign y17 = {(p6?p12:p8)};
endmodule
