module expression_00481(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd0)?(-2'sd1):(5'd27))?(5'd24):((4'sd0)?(3'd2):(-4'sd1)));
  localparam [4:0] p1 = (~((2'sd0)?(2'sd0):(3'd3)));
  localparam [5:0] p2 = (|(~(!{1{(-5'sd14)}})));
  localparam signed [3:0] p3 = ((((3'sd3)!=(4'sd4))|((2'd2)&&(4'd13)))>{1{{((4'd2)<(-3'sd0)),((4'd4)^~(3'sd2)),(5'd2 * (5'd4))}}});
  localparam signed [4:0] p4 = (2'd1);
  localparam signed [5:0] p5 = (-(4'sd0));
  localparam [3:0] p6 = ((!(4'd2))!==((2'd3)<<<(3'd5)));
  localparam [4:0] p7 = ((4'd8)^~(3'd5));
  localparam [5:0] p8 = ((-2'sd0)==(2'sd1));
  localparam signed [3:0] p9 = (2'sd1);
  localparam signed [4:0] p10 = (((3'sd3)?(-5'sd14):(5'd18))<<<((2'sd0)?(3'd6):(-5'sd9)));
  localparam signed [5:0] p11 = ((~&((~(3'sd0))>((-2'sd1)-(2'sd1))))>>>(((3'd2)>>(3'd1))+((2'd3)<<(-3'sd1))));
  localparam [3:0] p12 = (3'd4);
  localparam [4:0] p13 = (-(5'd29));
  localparam [5:0] p14 = (5'sd5);
  localparam signed [3:0] p15 = (^{2{{1{({2{(5'd16)}}^~((4'd9)!=(5'd30)))}}}});
  localparam signed [4:0] p16 = ((5'sd9)|(5'd17));
  localparam signed [5:0] p17 = (((5'sd2)&&(-(2'd0)))?((4'sd5)>>>(~(3'd4))):((2'd0)<(~&(5'd30))));

  assign y0 = (p3&&p1);
  assign y1 = (((p8%p15)?(p1?p5:p13):(p11>>p4))^~((~|(!p15))^(b1?p13:p14)));
  assign y2 = (~&(~|{3{(-5'sd6)}}));
  assign y3 = ({4{p3}}<(p2<p7));
  assign y4 = (~(3'd0));
  assign y5 = ((((|p6))==(3'd0))^(~&(&$signed({(p10-p9)}))));
  assign y6 = (({2{a5}}?{4{p11}}:(b2<=b4))?(2'd1):((a1==p2)?(p9&&b1):(b3!=a3)));
  assign y7 = ((b4<<<b0)||(-4'sd5));
  assign y8 = ((b0)>=(a1));
  assign y9 = (|(~|({(b5<<<p6),(p14?p9:b4),(|a2)}?$unsigned((b3?a0:b3)):$signed({3{b0}}))));
  assign y10 = (+(+(|($signed($signed($unsigned({b3,b5})))<{(b0),$unsigned(a3)}))));
  assign y11 = (p7&a4);
  assign y12 = ((p7-p9)>>>(-4'sd2));
  assign y13 = (4'd14);
  assign y14 = (~|(!$signed((~|($unsigned((|(|(p4!=p10))))=={(p15||p1),(~^p2)})))));
  assign y15 = $signed({{($signed($signed(a3))=={p5,b1,p15})}});
  assign y16 = (~^{(5'd16),(!(-4'sd0))});
  assign y17 = (($signed({p3,p0})^(((p14))))-((6'd2 * (p2>=p6))|$signed({p2,p11,p10})));
endmodule
