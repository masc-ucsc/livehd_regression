module expression_00345(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((5'd3)^~(-2'sd1))>=(5'd25))};
  localparam [4:0] p1 = {{2{(3'd0)}},((3'd5)!==(2'sd1))};
  localparam [5:0] p2 = (+(+((~^(-(~|(4'd12))))|(3'sd3))));
  localparam signed [3:0] p3 = (({2{(-3'sd2)}}<={3{(-2'sd0)}})<<{3{(-2'sd1)}});
  localparam signed [4:0] p4 = (&{1{(3'd7)}});
  localparam signed [5:0] p5 = ((((5'd0)<<(5'sd8))!==((5'd4)>>(2'd3)))&&(((5'd5)>>>(-3'sd2))<=((2'd2)&(-4'sd3))));
  localparam [3:0] p6 = (-(~^(~&(^(~&(~&(&(~|(~&(~&(|(!(~&(&(-3'sd2)))))))))))))));
  localparam [4:0] p7 = {(~(5'd8)),(+{((2'd0)<<(2'd3))})};
  localparam [5:0] p8 = ((-5'sd4)>(4'sd4));
  localparam signed [3:0] p9 = (({3{(2'd1)}}&{4{(5'd22)}})|(~^(~(!((&(3'd4))||(3'd4))))));
  localparam signed [4:0] p10 = ({1{(((-2'sd0)?(-2'sd1):(3'sd0))!=={4{(-5'sd14)}})}}&&{1{({4{(-5'sd7)}}^~{1{(2'sd0)}})}});
  localparam signed [5:0] p11 = (({1{((5'd7)&&(-4'sd4))}}|(~^((2'sd0)===(5'd19))))&({1{(-3'sd1)}}?(^(-4'sd1)):{2{(-3'sd2)}}));
  localparam [3:0] p12 = (((-2'sd1)||(4'd8))?((3'sd2)?(5'sd4):(4'sd4)):((5'd23)?(2'd0):(4'd0)));
  localparam [4:0] p13 = (+(~^(((~^{(4'd1),(3'd7)})&(5'd2 * (3'd5)))+(~&({(-5'sd5),(-3'sd3),(-3'sd1)}>>(-(2'd3)))))));
  localparam [5:0] p14 = (~&((((2'd2)^~(-5'sd3))+((2'd3)===(-2'sd0)))-(|(((3'sd0)<<(4'sd1))<<<(~^(-2'sd0))))));
  localparam signed [3:0] p15 = (|((6'd2 * ((4'd6)*(5'd2)))>=(((-3'sd0)<=(2'd2))<=((4'd6)<<(-2'sd1)))));
  localparam signed [4:0] p16 = (-4'sd6);
  localparam signed [5:0] p17 = ((2'd2)?(2'd0):(-5'sd9));

  assign y0 = (~^(~&({(p1<<<a3),(3'sd3),{a2,b2}}^~({b2,a5,b2}!==(~(5'd4))))));
  assign y1 = (&b2);
  assign y2 = ((((a5>>p0)>>>(a4<=b5))<=(+(~&(b2))))<<<(-((|(b0>=a5))===((b0^~a0)))));
  assign y3 = (^({4{b2}}!=(p16!=p6)));
  assign y4 = (3'sd1);
  assign y5 = {3{(({1{b1}}))}};
  assign y6 = ((b5?p13:p8)?((p2>>p14)<(p4?p0:b4)):((p12>>p6)*(p10?p9:p0)));
  assign y7 = {{(&(a4<=a1))},(^(b1<<p10))};
  assign y8 = {p6,p14,p7};
  assign y9 = {4{(+{4{b0}})}};
  assign y10 = (~&(-3'sd3));
  assign y11 = (+(~&(5'd14)));
  assign y12 = ((5'sd14)?(2'd2):((b0?b5:b5)>>(b1)));
  assign y13 = (-({2{p15}}+(a5<b2)));
  assign y14 = (b2<a3);
  assign y15 = {{({b1}|{a3,b1,b2}),({3{a1}}||{1{a2}}),{4{p16}}}};
  assign y16 = (5'd2 * (3'd1));
  assign y17 = (^{1{{1{(~p2)}}}});
endmodule
