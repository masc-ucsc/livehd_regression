module expression_00488(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'sd0)+(3'sd3))+(5'sd15))&&(-2'sd1));
  localparam [4:0] p1 = (|{1{(!(~^(4'd5)))}});
  localparam [5:0] p2 = (~^{2{(-4'sd3)}});
  localparam signed [3:0] p3 = (~&(-2'sd0));
  localparam signed [4:0] p4 = ((2'sd0)<(4'd3));
  localparam signed [5:0] p5 = ({4{(4'd11)}}<<<{1{{4{(4'd9)}}}});
  localparam [3:0] p6 = ({(-3'sd1),(4'sd6)}^{(-5'sd0),(-5'sd11),(5'sd13)});
  localparam [4:0] p7 = {{((5'd11)<=(3'd2))},{(-4'sd2),(4'd6)},{(3'd3),(3'd1),(-5'sd7)}};
  localparam [5:0] p8 = (((3'sd0)?(-5'sd8):(2'd0))<<((5'd25)?(4'd3):(-3'sd3)));
  localparam signed [3:0] p9 = (5'd18);
  localparam signed [4:0] p10 = ((((5'sd11)^~(2'd1))>>>((2'sd0)?(3'sd3):(-4'sd7)))+(((3'd0)?(4'd4):(5'sd7))|(4'sd6)));
  localparam signed [5:0] p11 = {({(2'd1),(5'sd14)}?{1{(4'd13)}}:{(3'd7),(2'd1)}),{{(2'sd1),(2'd1),(-3'sd2)},{2{(5'sd12)}},((5'd30)>>(2'sd0))}};
  localparam [3:0] p12 = (((4'sd0)?(-2'sd0):(3'd2))=={((2'd0)<=(3'd3)),((-2'sd1)?(4'd9):(5'sd5))});
  localparam [4:0] p13 = (+(2'd3));
  localparam [5:0] p14 = (~^(~&(-5'sd14)));
  localparam signed [3:0] p15 = (^(+((5'd2 * (4'd10))/(3'sd0))));
  localparam signed [4:0] p16 = (~^((3'sd3)===(((2'd1)&&(4'd2))+((4'sd3)!==(5'd18)))));
  localparam signed [5:0] p17 = (~((((-2'sd1)?(3'sd1):(-4'sd4))?(5'sd5):((4'd15)==(4'sd1)))||((5'sd1)?((4'd5)<<<(4'd8)):(-5'sd8))));

  assign y0 = ($signed((4'd8))?(~&(!$signed(b4))):(4'd5));
  assign y1 = {(!(p0?p0:p15)),(b0==p1),(-{1{p2}})};
  assign y2 = ({4{a4}}>>(~^a1));
  assign y3 = {2{(|((^p5)?(b2+b2):(|a3)))}};
  assign y4 = (5'd23);
  assign y5 = {(p6>p15),{p13,p14}};
  assign y6 = ((b2>>>a5)<=(a1-a4));
  assign y7 = ((a3>>>a4)?(b5?b2:b1):(a5<=b0));
  assign y8 = (4'd7);
  assign y9 = {{(b0?p17:p8),(b2?a3:p3),(p5?p12:p15)},{(a3?p7:b3),(b2===a4)}};
  assign y10 = (5'd24);
  assign y11 = ({(p12<a1),(a1^a5)}?({b0,b1}>=(a1^p8)):{1{(6'd2 * {a2,b1})}});
  assign y12 = {({a4}>>>(b1||a2)),((b2!==b3)!==(b4>b2)),(-(~|(~|$signed(a3))))};
  assign y13 = {1{({3{{1{b2}}}}?(6'd2 * {(4'd15)}):((b2|a2)^(3'sd0)))}};
  assign y14 = $unsigned((((b0))*(b2<<<b2)));
  assign y15 = ((~((b5-b3)?(~p11):(a5<<<a1)))==(^(+(a3?a3:a0))));
  assign y16 = ({4{(a0<b4)}}||$unsigned(($signed(({4{b3}}>(a2==b1))))));
  assign y17 = {2{(~|p1)}};
endmodule
