module expression_00171(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{(4'd11)}}+{(2'd2),(4'sd7),(-5'sd0)});
  localparam [4:0] p1 = (2'd0);
  localparam [5:0] p2 = ((3'sd0)?(5'd24):(2'sd0));
  localparam signed [3:0] p3 = (~&{(+((3'sd0)?(3'sd3):(-4'sd0))),((4'd12)?(2'd0):(3'd7)),(+(2'sd0))});
  localparam signed [4:0] p4 = {2{(-2'sd1)}};
  localparam signed [5:0] p5 = (((5'sd10)/(3'd4))!=(2'sd1));
  localparam [3:0] p6 = (~^(-(&(&{4{(4'd9)}}))));
  localparam [4:0] p7 = ((~^{(((4'sd7)?(2'd3):(4'd5))?(-(5'd26)):{(-5'sd2)})})!=(~|((~^((2'sd0)<<<(3'd3)))+((2'sd1)>>>(5'd21)))));
  localparam [5:0] p8 = (4'd2 * (3'd0));
  localparam signed [3:0] p9 = {((((-5'sd4)?(5'd28):(2'sd1))==((5'd9)^~(-4'sd1)))>(((3'sd0)?(5'sd2):(4'd4))?((5'd10)|(4'sd0)):{(3'sd0),(-4'sd7)}))};
  localparam signed [4:0] p10 = (((3'sd0)?(4'd7):(5'd13))?((3'd5)?(3'd3):(2'd1)):((5'sd2)?(2'd3):(2'd1)));
  localparam signed [5:0] p11 = {1{(-5'sd13)}};
  localparam [3:0] p12 = {(4'd5),(3'd6)};
  localparam [4:0] p13 = ((3'd1)!=(((5'sd13)===(5'd19))!=((-5'sd11)<=(5'd17))));
  localparam [5:0] p14 = (~&((~^(~^(!(+(5'd2 * (2'd0))))))|(~&(|{{(4'd12)},((2'd3)-(-5'sd1))}))));
  localparam signed [3:0] p15 = (((4'd1)>>>(3'd0))&((4'sd0)?(-5'sd10):(4'd12)));
  localparam signed [4:0] p16 = (((4'sd6)&(-5'sd0))!==((-3'sd0)?(5'd29):(-3'sd0)));
  localparam signed [5:0] p17 = (((5'd22)?(2'd1):(-5'sd4))!=(3'sd1));

  assign y0 = ((~|((+(((~^p0)>=(p1&b3))))-((&(~|$unsigned((p6<<<p15))))))));
  assign y1 = (~|(2'd1));
  assign y2 = (((|(p12))>>>$signed((a0>=p17)))<$unsigned(((a5<<p16)<=(+a5))));
  assign y3 = ((a1<p14)>(b4<=b1));
  assign y4 = (({a1,b1}===(a1&b5))!={(b3>=b1),(5'd2 * p13),(4'd2 * b0)});
  assign y5 = $unsigned(((($unsigned({$signed((^(3'sd3))),$signed((+(|p6))),({{p13,p7,p8}})})))));
  assign y6 = (&((6'd2 * p8)>($signed(b0))));
  assign y7 = (&({(p17<p2),(p9^p5)}|((p14>=p8)^(-{3{p2}}))));
  assign y8 = ({1{((|(-p10))-(b4||a2))}}^{1{((b1<b2)?{3{p2}}:(-3'sd0))}});
  assign y9 = (-5'sd11);
  assign y10 = ((((a0<a0)|{2{a1}})<=$unsigned((p13<<b4)))<<<(!(&(~^((b3<b4)>>(b4>>>b1))))));
  assign y11 = {((p15?b4:p16)?(b4?a1:p8):(a3&&a2)),({4{b3}}?{4{a4}}:(^{p2,a1}))};
  assign y12 = (|(~((5'sd15)?(p0<<p13):(a1?p0:p8))));
  assign y13 = ({4{{3{b2}}}}^~((^(~^(~|{4{p12}})))<<<((~b3)||(a5<=p5))));
  assign y14 = ({{(-3'sd2)}}<{{{p13,p7,b0}}});
  assign y15 = ($signed((!(3'd7)))^$signed((|$unsigned(b3))));
  assign y16 = (-(~^(~(b2?a3:b2))));
  assign y17 = (((b3&p11)?(p1+a5):(p10&&p17))!=({2{{1{a1}}}}+{1{((b5^~b2)<<(b4===a0))}}));
endmodule
