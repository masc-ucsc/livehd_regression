module expression_00466(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((((-3'sd3)&(4'd14))>=((4'sd5)/(-5'sd3)))+(((-3'sd1)<<<(2'd2))<=((5'd11)!=(3'd2))))^~((((5'sd14)>=(2'd2))!==((5'sd1)||(5'd12)))+(((-3'sd1)>>>(3'd5))!=((2'd1)>=(3'd3)))));
  localparam [4:0] p1 = ((((-5'sd13)<<<(2'd0))>((3'sd1)||(2'd1)))^(((5'd21)?(-5'sd0):(2'd0))<<{1{((-5'sd13)>=(4'sd4))}}));
  localparam [5:0] p2 = (^{((-3'sd1)!={(-3'sd0),(-3'sd1),(-3'sd0)})});
  localparam signed [3:0] p3 = (~&(&((((-2'sd0)?(-5'sd12):(-3'sd0))!==(5'd2 * (3'd0)))>=((~&(4'd13))<(5'd2 * (3'd6))))));
  localparam signed [4:0] p4 = (-4'sd4);
  localparam signed [5:0] p5 = (((~(2'd0))/(3'sd0))>>(5'd29));
  localparam [3:0] p6 = (~&((4'd3)&&(4'd12)));
  localparam [4:0] p7 = {4{{4{(5'sd4)}}}};
  localparam [5:0] p8 = ((~^(!((-3'sd3)?(3'd1):(2'd2))))?{2{(2'd0)}}:((5'd16)?((4'd14)?(-2'sd1):(3'sd2)):(|(-3'sd0))));
  localparam signed [3:0] p9 = {2{((5'd4)&&((-4'sd4)===(3'd6)))}};
  localparam signed [4:0] p10 = (~^(~^((4'd13)?(3'sd3):(-4'sd2))));
  localparam signed [5:0] p11 = (~(5'd2 * (|(^(3'd7)))));
  localparam [3:0] p12 = (((5'd27)!==(2'd0))>((3'd3)|(5'd1)));
  localparam [4:0] p13 = ((((5'sd4)?(2'sd1):(-5'sd5))?(~^(4'd4)):((4'sd2)?(2'd0):(-2'sd0)))?((+(-4'sd1))^(~(5'd5))):(&((-(2'd1))/(2'd1))));
  localparam [5:0] p14 = ((((3'd2)-(4'sd0))<<((3'sd2)^~(5'd10)))<<{((4'd4)<<(-4'sd7)),{2{(-5'sd14)}}});
  localparam signed [3:0] p15 = {2{(&(^{3{(2'd2)}}))}};
  localparam signed [4:0] p16 = (&(((!(5'd26))===((-5'sd11)?(-3'sd1):(4'd13)))?(((2'd2)-(5'd9))+((-3'sd0)^(3'd4))):(((2'sd0)^(-5'sd9))-((5'd9)?(2'd0):(4'd11)))));
  localparam signed [5:0] p17 = ((|({(5'sd8),(-4'sd2)}&((4'd14)<=(3'd5))))>>{(~&(3'd0)),((3'd3)<<(2'd2)),{(4'd15)}});

  assign y0 = ((p12+p5)?(a4<=p6):{1{(!a3)}});
  assign y1 = (+(((($unsigned((~|$unsigned((^(+$signed((b2))))))))))));
  assign y2 = ((b0===a2)?(&(p7<<p4)):(p8?p8:b1));
  assign y3 = $signed($unsigned($unsigned({$signed({1{{p12,p5}}}),$signed(({4{p13}})),{{p2},{p5,p0}}})));
  assign y4 = {{{{((-p8)==(p7?p17:a5))},((p3?p3:p15)|(b2?p12:a2)),({a5,p8}?{p2}:(p9?b3:b2))}}};
  assign y5 = (4'd1);
  assign y6 = (4'sd3);
  assign y7 = (a0?b0:b2);
  assign y8 = (~&{$signed({a2,p2,b1}),((a5?b1:b0)),(a5-a5)});
  assign y9 = (3'd0);
  assign y10 = (3'sd0);
  assign y11 = ({(5'd10),{2{p5}},{p15}}?(3'd7):(3'd4));
  assign y12 = {1{(&(~{3{(a0)}}))}};
  assign y13 = (^{2{(p3<<<p10)}});
  assign y14 = ({{b4,p7},(^b1),(a2?b2:b0)}?(+(&(b5!=a3))):{2{(p1?p0:a5)}});
  assign y15 = (|{1{(({3{{2{p14}}}}+{1{(-{2{{1{b4}}}})}}))}});
  assign y16 = ((~^{{{b1,b2}}})<(4'd2 * {p1,a2,a1}));
  assign y17 = (4'sd4);
endmodule
