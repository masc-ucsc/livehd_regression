module expression_00972(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'sd9)>=(4'd1))<{3{(-3'sd3)}});
  localparam [4:0] p1 = ((-{1{(3'sd3)}})?((2'd3)?(4'd8):(2'd2)):((3'sd3)^(5'd9)));
  localparam [5:0] p2 = (|(5'd29));
  localparam signed [3:0] p3 = (((-4'sd7)^(4'd9))<<{(2'd0),(3'sd3),(4'd4)});
  localparam signed [4:0] p4 = (+{(^{({(-2'sd0)}===((2'd2)>>>(5'd0)))})});
  localparam signed [5:0] p5 = ((-5'sd13)?(-5'sd13):(4'd9));
  localparam [3:0] p6 = {(-2'sd1),(|((-5'sd15)&(3'd5)))};
  localparam [4:0] p7 = (2'd2);
  localparam [5:0] p8 = (~|((2'd3)<=(4'sd4)));
  localparam signed [3:0] p9 = {1{(4'd11)}};
  localparam signed [4:0] p10 = (~|(5'd2 * (5'd11)));
  localparam signed [5:0] p11 = (({(4'd2),(-5'sd12),(5'sd1)}!=((-5'sd2)?(-3'sd0):(5'sd10)))?{(5'd15),(4'd14),(4'sd5)}:(2'd1));
  localparam [3:0] p12 = ((((5'd25)||(2'sd0))?((4'sd0)?(-4'sd3):(5'd17)):{2{(4'd10)}})+{4{((5'd14)==(2'sd0))}});
  localparam [4:0] p13 = {(2'd2)};
  localparam [5:0] p14 = ((((-5'sd8)>>(2'd1))||((-5'sd15)?(5'd1):(3'd6)))+(~&((~|(4'sd4))?(~(-3'sd1)):(~^(-5'sd11)))));
  localparam signed [3:0] p15 = ((-(-(-3'sd1)))|(+(((4'd13)^(3'd0))^((5'd30)>>>(3'd2)))));
  localparam signed [4:0] p16 = ((~&(+{2{{1{(~&(3'd6))}}}}))<<<(-{2{((5'sd11)===(2'sd1))}}));
  localparam signed [5:0] p17 = ((((3'd4)?(3'd2):(4'sd2))<<<(((4'd7)-(4'd14))&&((4'd5)?(-2'sd0):(4'd6))))^~((+((2'sd0)+(3'd0)))||(~|(-((2'sd0)===(4'd7))))));

  assign y0 = {1{(a1>a0)}};
  assign y1 = ((p4<<<b4)?{a4,a1}:{a3,p17});
  assign y2 = (~(~&(+({1{(b5===a4)}}===(~^{2{a1}})))));
  assign y3 = (+(~|$unsigned((5'd18))));
  assign y4 = (((a4<b2)^(a5>=b2))?((a4!==a3)&&(a0?a0:p11)):((a1+p10)>=(a1<=b5)));
  assign y5 = {({((p10<<b4)),{p6,b2,a0},(~^{a2,b5,a4})})};
  assign y6 = (5'sd7);
  assign y7 = (b1<a5);
  assign y8 = (3'd0);
  assign y9 = {a1,p8};
  assign y10 = ({1{a4}}||{3{a1}});
  assign y11 = (|({$unsigned({p6,p9,a4})}||({b3}||(b5!==b5))));
  assign y12 = (!$signed((|$signed($unsigned((^((~^(^((|(^p7))))))))))));
  assign y13 = (5'sd11);
  assign y14 = ((~^({1{(b1>b3)}}&&(a2===a2)))|{4{(3'sd3)}});
  assign y15 = ((+((b3|p15)<(+(~^b1))))>=((&{a3})>>>{{p15,p3,p2}}));
  assign y16 = $signed((p0>>p1));
  assign y17 = {2{(~p1)}};
endmodule
