module expression_00809(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((4'd1)^~(2'd2))};
  localparam [4:0] p1 = ((3'sd2)-{{{(5'd10)},((2'd3)?(2'd3):(-4'sd3))}});
  localparam [5:0] p2 = ({2{{3{(-4'sd7)}}}}||(~|((2'sd1)?(3'sd1):(2'd2))));
  localparam signed [3:0] p3 = (5'd26);
  localparam signed [4:0] p4 = (((4'd6)===(-5'sd13))?(~^(~&(-2'sd1))):(-5'sd4));
  localparam signed [5:0] p5 = ((4'd2 * (3'd7))-((4'd5)?(-5'sd11):(4'd5)));
  localparam [3:0] p6 = ((3'd1)?(~(-{3{(3'sd3)}})):(((3'd6)?(3'sd2):(5'd25))^~((2'd2)?(-5'sd3):(4'sd7))));
  localparam [4:0] p7 = {3{{(-5'sd4),(2'sd1),(5'd18)}}};
  localparam [5:0] p8 = {2{(+(+{1{((4'sd1)>(-4'sd1))}}))}};
  localparam signed [3:0] p9 = (((3'sd2)>>>(4'd14))<(6'd2 * (5'd15)));
  localparam signed [4:0] p10 = (^(((5'd23)%(4'd0))^((-2'sd1)!==(-4'sd0))));
  localparam signed [5:0] p11 = ((((4'd9)<<(4'sd5))?((2'sd0)?(2'd0):(4'd15)):((3'd4)>>>(3'd3)))>>>({4{(5'd16)}}?((3'd4)?(-3'sd2):(5'sd8)):{1{(4'sd4)}}));
  localparam [3:0] p12 = (((!(4'd2))<<(&(5'd1)))^~{4{(3'd7)}});
  localparam [4:0] p13 = (&({(2'd3),(4'sd4),(3'sd0)}<<<(&(~|(6'd2 * (3'd0))))));
  localparam [5:0] p14 = {({{3{(5'sd11)}},{3{(4'sd7)}}}==(5'd2 * (&{(2'd1),(5'd9),(2'd2)})))};
  localparam signed [3:0] p15 = (~^(+(^({(~(-3'sd0)),{(-5'sd12),(2'd3)}}^((2'sd1)^{3{(4'd1)}})))));
  localparam signed [4:0] p16 = (|(~|(3'd6)));
  localparam signed [5:0] p17 = (~^({(+(4'sd1)),{(2'd3)},(4'd2)}<<(4'd1)));

  assign y0 = (5'd2 * {a0,a1});
  assign y1 = ((+p13)?(~|p4):{3{p7}});
  assign y2 = ((((|(p11<p6)))<<<({3{a5}}>>>(b4^b5)))==(((b2>>>b3)>>>(b2>>p17))));
  assign y3 = (((b4===a3)+(p14&&b2))&&((~&(p6<<p6))>>(b1||p1)));
  assign y4 = (~&(-4'sd0));
  assign y5 = (-3'sd1);
  assign y6 = ((5'sd13)^{(-2'sd1),(a4!==a2)});
  assign y7 = {1{{1{(+((a4)?(a3):$signed(p2)))}}}};
  assign y8 = ((a5===a0)<<<{3{a1}});
  assign y9 = (~^{(!{(-2'sd1),(^((~^a3)=={a1})),{(~^p10),(|a5),(+b3)}})});
  assign y10 = ((a0!==a5)>{p7,p4});
  assign y11 = ((^((p0?a4:p5)<<<(p6||p6)))+(+(~|(b5?b2:a2))));
  assign y12 = (+{4{((p3<p3)>>>(~&p10))}});
  assign y13 = $signed(((2'd2)));
  assign y14 = ((^(&(a3^~p15)))&((5'd2 * p7)^(|a0)));
  assign y15 = (!(&(!(&(!(~^(~(~&(-(&(|(~^(-(~^(^p11)))))))))))))));
  assign y16 = ((((a2===a2)===(b4>>b4))<<((b5-a5)>=(5'd2 * a1)))|((a3-a2)/a1));
  assign y17 = (!(~$signed(((^(~^(~(~(p17)))))<<({a1,a3,b2}!=(&(-b1)))))));
endmodule
