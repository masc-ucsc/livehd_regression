module expression_00679(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-2'sd0)?(3'sd0):(2'sd1));
  localparam [4:0] p1 = ((4'd2)>={{((-5'sd6)?(4'sd1):(-2'sd0))}});
  localparam [5:0] p2 = ((~(5'd22))?((-5'sd9)?(4'd2):(3'sd0)):((5'd11)?(2'd0):(-2'sd0)));
  localparam signed [3:0] p3 = (^(~^{(+(^(4'sd0))),(~|{(-5'sd13),(3'd0),(5'd16)})}));
  localparam signed [4:0] p4 = (!{{(-4'sd3),(3'd4)},(~{(5'd14),(2'd3)})});
  localparam signed [5:0] p5 = (((3'd6)^(2'd1))<=((5'sd3)<<(2'd3)));
  localparam [3:0] p6 = (((2'd1)>=(-5'sd10))<((2'd3)==(3'd3)));
  localparam [4:0] p7 = {(((5'd13)>>(-3'sd3))?{(3'd1),(2'd1),(4'd14)}:((-2'sd0)>>(2'sd0))),(((4'd14)?(-5'sd6):(-4'sd6))?((3'd6)?(-5'sd6):(3'd6)):((2'd0)^~(2'd3))),({4{(2'd3)}}+{(4'd3),(-2'sd0),(-3'sd1)})};
  localparam [5:0] p8 = (({(3'd1),(-3'sd2)}>>>((2'd1)|(4'd10)))!==(((-2'sd1)^~(4'd15))^~(^(5'd13))));
  localparam signed [3:0] p9 = (~(~^((~|(((3'd7)||(3'd7))-(~^(^(5'd13)))))<<(!((+(|(2'd2)))!=(-((5'd8)<=(3'sd0))))))));
  localparam signed [4:0] p10 = {3{(((5'd7)>>>(2'sd1))^~(5'd2 * (2'd3)))}};
  localparam signed [5:0] p11 = {{(((2'd0)>>(4'd11))>>((3'sd1)===(5'd9)))},(((-3'sd2)!==(4'd7))+((3'd4)!=(-2'sd1)))};
  localparam [3:0] p12 = ((4'd3)/(4'sd1));
  localparam [4:0] p13 = ((((3'd5)?(-3'sd0):(3'sd3))?((4'sd3)||(5'd31)):((-2'sd1)+(4'sd5)))<=(|(~|((5'd2 * (4'd1))|(-3'sd0)))));
  localparam [5:0] p14 = (|(5'd2 * ((4'd4)<<<(5'd23))));
  localparam signed [3:0] p15 = (((3'd0)>(2'd0))?(4'd12):{(5'd30),(2'sd0),(5'sd7)});
  localparam signed [4:0] p16 = (4'd1);
  localparam signed [5:0] p17 = {({3{(2'sd1)}}?(^(5'd12)):{(2'sd1),(-4'sd7),(-2'sd1)}),{{(-3'sd3),(5'sd10)},((5'd11)!==(4'sd0))}};

  assign y0 = {4{(~{4{a0}})}};
  assign y1 = (-2'sd1);
  assign y2 = ({{{(p6!=b0),{a3,a3,p11}}}}>>>({1{{p8,p7}}}<={4{p16}}));
  assign y3 = (~(-2'sd1));
  assign y4 = (((-(-(b2-a2)))&&((a4<p14)|(b5<<b2)))<((b2!=a3)/b5));
  assign y5 = ((~^(a2==p1))!={p11,a5,b2});
  assign y6 = {3{(5'd19)}};
  assign y7 = (((p3<p12)?(b1&&b2):{2{b5}})!={2{((a2?a1:b4)>={4{a4}})}});
  assign y8 = (((p11?p5:b2)?(2'd1):(a1?a0:p2))?{3{{4{p15}}}}:((p16>b2)?{1{a4}}:(a0?a3:b4)));
  assign y9 = {1{((p3?b5:a0)|(+(a0>>>b1)))}};
  assign y10 = {((!a4)?{a3}:{p10}),{(~(&b4)),{b2,p5}},(+({b3,a5,a3}+(a1^~b2)))};
  assign y11 = (5'd15);
  assign y12 = {4{{p7,p16}}};
  assign y13 = {$signed(p10),{b2},{p6,p2,a3}};
  assign y14 = ({2{(p15?p6:a0)}}|{2{(-4'sd4)}});
  assign y15 = (+((b4^~p0)-{2{p17}}));
  assign y16 = (2'd3);
  assign y17 = (+((-((p11^p15)^~(b0^~a2)))>=(!((5'd2 * p12)%b1))));
endmodule
