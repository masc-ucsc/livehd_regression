module expression_00836(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~^(4'sd5))?(^(-2'sd1)):((-3'sd0)?(-5'sd12):(3'sd1)))==={4{(3'd1)}});
  localparam [4:0] p1 = ({(-3'sd1),((2'd3)|(5'd10))}!={{((3'sd2)&(5'sd13))},(&(~|(3'sd0)))});
  localparam [5:0] p2 = {3{{4{(-4'sd6)}}}};
  localparam signed [3:0] p3 = (4'sd2);
  localparam signed [4:0] p4 = ((3'sd2)&(5'sd5));
  localparam signed [5:0] p5 = ({1{{3{(4'd4)}}}}!==(((3'd1)?(4'sd2):(5'd2))?((-5'sd5)==(2'd3)):((4'd5)?(4'd0):(3'sd0))));
  localparam [3:0] p6 = (^(~&(((2'd3)/(-4'sd6))+(&(~&(-4'sd6))))));
  localparam [4:0] p7 = {(-4'sd6),((4'd9)<<{(5'sd9),(-3'sd3),(5'sd13)})};
  localparam [5:0] p8 = ((((2'd2)?(5'd9):(-2'sd0))!==((4'd14)?(5'sd10):(4'd0)))<<{1{((3'sd1)?(5'sd4):(4'd7))}});
  localparam signed [3:0] p9 = (((-4'sd7)>=(-4'sd6))==(4'd2 * (4'd7)));
  localparam signed [4:0] p10 = ({1{{1{((2'd3)<{2{(5'sd5)}})}}}}!=((((5'd4)||(-5'sd3))==(3'd2))^~(3'sd1)));
  localparam signed [5:0] p11 = (-5'sd7);
  localparam [3:0] p12 = (((3'd4)?(~(~|(3'd5))):(-(3'd3)))|(3'sd3));
  localparam [4:0] p13 = (!{3{{(-3'sd1),(-5'sd6)}}});
  localparam [5:0] p14 = {3{(5'd6)}};
  localparam signed [3:0] p15 = ((((2'sd0)>>>(2'd3))!==((2'sd0)+(3'd2)))==(((3'd0)>(4'd1))/(4'sd0)));
  localparam signed [4:0] p16 = (&(2'sd1));
  localparam signed [5:0] p17 = {4{(+{3{(2'd3)}})}};

  assign y0 = $signed({3{(^b4)}});
  assign y1 = (^(-(((-(p1^~p16))||(~|(~&p10)))+($unsigned((~^p2))<=(p3|a1)))));
  assign y2 = ((-3'sd1)||{4{p3}});
  assign y3 = ($signed(a1)?(b3<<<p10):{2{b1}});
  assign y4 = ({(~|(!(~&$unsigned({p9,p5,p5})))),(+(|((~|(~{p4})))))});
  assign y5 = ((~(((&b4)!=(p1+b0))!=((p9*a4)%b3)))!=(^((!(b4||a3))&&(!(b0+p8)))));
  assign y6 = {4{{4{b2}}}};
  assign y7 = {$signed(b1),{p13,b3},(b1)};
  assign y8 = (~((4'd11)));
  assign y9 = ({a5,p5}?{4{b4}}:(a2?p1:a0));
  assign y10 = (((2'd2))<<<((5'sd10)^(-3'sd1)));
  assign y11 = (^{2{{3{$signed($unsigned(p12))}}}});
  assign y12 = {2{{1{(2'sd1)}}}};
  assign y13 = {$unsigned((p10)),$signed((p4?p12:p17)),(~^(!p7))};
  assign y14 = {1{(-3'sd3)}};
  assign y15 = (((p12?p7:p2)==(p13>=p0))?({p3,p3,p17}?(p14||p8):(p1?p17:p7)):((p4<<p3)?(2'd1):(p11||p9)));
  assign y16 = (((a1?p2:p4)%p0)>>>(p14?p12:p17));
  assign y17 = (2'd1);
endmodule
