module expression_00951(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+(~&(5'd4)))?((5'd28)?(2'd2):(4'd15)):((-5'sd8)?(4'd11):(4'd12)));
  localparam [4:0] p1 = (~^(((!(4'sd6))?(!(5'sd6)):((-4'sd3)<(-3'sd3)))<{4{(-2'sd0)}}));
  localparam [5:0] p2 = (5'd18);
  localparam signed [3:0] p3 = (&{{(2'd0),(5'd1),(4'sd0)},((!(-4'sd3))!=((5'd30)+(-3'sd3))),(4'd11)});
  localparam signed [4:0] p4 = (((-3'sd3)|(-5'sd3))+((-2'sd1)|(4'd1)));
  localparam signed [5:0] p5 = (^(~^(^(~|(|(&(-3'sd2)))))));
  localparam [3:0] p6 = ((+((2'd2)?(5'sd14):(-3'sd0)))^{4{(5'd12)}});
  localparam [4:0] p7 = {2{((+((4'd1)!==(4'd1)))<=((-4'sd0)>(4'sd5)))}};
  localparam [5:0] p8 = ({((5'd21)-(3'd2)),{(-5'sd2)},{(2'd3)}}>=({(4'd4),(-5'sd5),(3'd5)}^~((-2'sd1)!=(3'sd2))));
  localparam signed [3:0] p9 = (~&(~&(((^(5'd27))>((-2'sd0)<<<(2'd3)))<<(~(((3'd6)>(2'd0))>((5'd24)/(5'sd15)))))));
  localparam signed [4:0] p10 = {(~|(3'd2))};
  localparam signed [5:0] p11 = (^(~|(-(6'd2 * (!(~(4'd8)))))));
  localparam [3:0] p12 = ((~&(!{(5'sd2),(3'sd2),(2'd2)}))===({(-4'sd5),(3'd0)}!==(|((3'd2)&(-5'sd8)))));
  localparam [4:0] p13 = (-(-2'sd0));
  localparam [5:0] p14 = (~^(-(((-4'sd1)+(-5'sd3))>>>{(4'd9),(-5'sd14),(4'sd2)})));
  localparam signed [3:0] p15 = (+(4'sd7));
  localparam signed [4:0] p16 = ((5'd1)/(4'd15));
  localparam signed [5:0] p17 = (5'd13);

  assign y0 = ((~|(p10==p6))?(2'd1):(2'd3));
  assign y1 = {2{(p1?b4:p10)}};
  assign y2 = ((((b0-b3)%b5)&((b1*b2)>(a5/b2)))==(((p12==b2)!=(p4&b5))>>>((b0*a5)>>>(a3/a5))));
  assign y3 = (((-5'sd4)>>>{3{b1}})==={{3{(b1==a4)}}});
  assign y4 = (!p2);
  assign y5 = $signed((!$signed(({2{($unsigned((!((2'd0)||(2'd1)))))}}))));
  assign y6 = ((5'sd11)?((b3>>>b4)>=(b4?p5:a1)):(-(a3?p10:p7)));
  assign y7 = ((~(~|(p17?p12:p7)))?(^(^(p1?p10:p15))):(((p16?p9:p3)?(!p10):(p13))));
  assign y8 = ((p9?p7:b2)||(p16-p10));
  assign y9 = (3'd0);
  assign y10 = {1{(3'd5)}};
  assign y11 = (p9&&p1);
  assign y12 = (a2>a3);
  assign y13 = ({a0,b3}>={p2,p10,p8});
  assign y14 = ((b1&p11)?{(b5|a4)}:{4{b3}});
  assign y15 = {3{(&(&(5'sd2)))}};
  assign y16 = (5'd3);
  assign y17 = (!(({4{a1}}?(~^p5):(^b1))?({2{p15}}?(a5|p12):(p17>>>p0)):(~{2{(a5&p4)}})));
endmodule
