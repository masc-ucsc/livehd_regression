module expression_00305(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|(3'd3));
  localparam [4:0] p1 = (+{1{((|((-5'sd7)==(5'sd1)))-{1{((-3'sd0)?(4'd4):(4'd4))}})}});
  localparam [5:0] p2 = (((-3'sd3)?(4'd0):(5'd28))+{(5'd24),(4'd1)});
  localparam signed [3:0] p3 = (+(((5'd2 * (2'd1))>>>((2'sd0)&&(5'sd14)))>={(5'sd12),((4'd6)||(2'd3)),(2'd1)}));
  localparam signed [4:0] p4 = (((3'sd3)&(5'd7))!=((5'd18)>=(5'd5)));
  localparam signed [5:0] p5 = (!((&(3'sd2))?{1{(4'sd3)}}:((2'd3)<<<(3'd0))));
  localparam [3:0] p6 = (3'd6);
  localparam [4:0] p7 = {(|(~&(((^(4'd1))^{(-5'sd5),(4'd10)})&&((5'd21)^(3'sd2)))))};
  localparam [5:0] p8 = ((2'd1)>>(|{2{(2'd1)}}));
  localparam signed [3:0] p9 = (((3'sd1)!=(4'd3))+((3'sd3)&(4'd1)));
  localparam signed [4:0] p10 = ((~&(5'd5))>(2'd0));
  localparam signed [5:0] p11 = (&(((-5'sd7)^(-3'sd2))|((3'sd2)>=(2'd0))));
  localparam [3:0] p12 = (3'd2);
  localparam [4:0] p13 = {(2'd1),(3'sd1)};
  localparam [5:0] p14 = (~&((~|((~&(-3'sd1))>(+(2'd1))))===((|(-4'sd1))^~(+(-2'sd1)))));
  localparam signed [3:0] p15 = {4{{4{(2'd3)}}}};
  localparam signed [4:0] p16 = (~^(&(|(&(&(~&(~|(+(+(!(!((2'd2)?(5'd8):(2'd3)))))))))))));
  localparam signed [5:0] p17 = (((2'd2)?(4'd10):(3'd3))?(|(&(5'd0))):(~&((3'd6)?(-5'sd5):(-5'sd8))));

  assign y0 = (~^({1{(^{2{b0}})}}!=={3{(a1-b5)}}));
  assign y1 = (~(&((a2?b0:b4)<<<(a2?p11:b4))));
  assign y2 = ({(-4'sd5)}>={(b3<=a1),(b4>=a3)});
  assign y3 = (5'sd15);
  assign y4 = ((&(2'd0))<(4'sd7));
  assign y5 = (~&(~(+(-5'sd5))));
  assign y6 = (((&b0)?(b1):$signed(a3))?({p14,a3}?{p1,p3,p5}:$unsigned(a1)):(~|((a3?a0:p8)<=(~^(a1)))));
  assign y7 = ({1{{(p6|p13),(2'sd1)}}}>=((p2&p3)==(p8!=p10)));
  assign y8 = (-{((~(&(2'd2)))<={2{(p17|a2)}}),(+({(~^(-4'sd3))}>={2{{b3,p11,p11}}}))});
  assign y9 = (~^$unsigned((^((~^$signed(p1))?$signed((b0?p8:p5)):(~^(~^p3))))));
  assign y10 = (&{3{p16}});
  assign y11 = ({4{p13}}?$unsigned($signed((4'd9))):$signed({2{a1}}));
  assign y12 = ((~(+$signed($signed({1{(5'sd5)}}))))>>(5'sd3));
  assign y13 = ((a5>>a0)!==(a5));
  assign y14 = ((3'd2)^$signed({4{p0}}));
  assign y15 = ((((!(~^{2{a0}}))>=((a1?p17:b4)))));
  assign y16 = (-(((4'd13)==((a0>>>a4)|(a5>b4)))!=((-5'sd2)&&(5'd27))));
  assign y17 = {{(p8?b2:a4),(3'd2),{b5,b0}},({p11,a3}?(a0?a2:p12):{p6,p9,a5})};
endmodule
