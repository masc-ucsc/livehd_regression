module expression_00877(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'sd4)&(-5'sd9));
  localparam [4:0] p1 = {3{({2{(3'd6)}}==={3{(3'd6)}})}};
  localparam [5:0] p2 = ((-3'sd1)<<<({1{{(3'd2)}}}>(3'sd1)));
  localparam signed [3:0] p3 = ((~^(((-3'sd2)?(-2'sd1):(4'd3))?{2{(4'd3)}}:((-2'sd0)!=(4'd13))))&(((5'd22)||(2'sd0))^~(-{3{(2'd3)}})));
  localparam signed [4:0] p4 = (+((-2'sd1)>=(2'sd0)));
  localparam signed [5:0] p5 = ({1{(4'd12)}}+((3'sd0)!==(-5'sd15)));
  localparam [3:0] p6 = {2{(3'sd2)}};
  localparam [4:0] p7 = {(+{((!(-2'sd1))+{2{(-2'sd1)}}),((5'd12)?(4'sd5):(2'd0)),(-((4'sd4)>>(5'd28)))})};
  localparam [5:0] p8 = (-5'sd11);
  localparam signed [3:0] p9 = (-4'sd0);
  localparam signed [4:0] p10 = (3'd2);
  localparam signed [5:0] p11 = (~|{(-{1{{1{(|((((3'd3)|(3'd3))<((5'd4)<<(-3'sd3)))&{(+(2'd0)),((-2'sd0)<=(-4'sd0))}))}}}})});
  localparam [3:0] p12 = (((2'd2)^~(4'd7))?{(-5'sd6),(5'sd12),(3'sd0)}:((-5'sd5)&&(2'd0)));
  localparam [4:0] p13 = ((5'sd2)<<(5'd30));
  localparam [5:0] p14 = ((-5'sd6)*(-3'sd3));
  localparam signed [3:0] p15 = ((((4'd12)!=(4'd12))|(5'sd5))!==((2'sd0)>(2'd1)));
  localparam signed [4:0] p16 = (&((3'd2)<<(2'sd1)));
  localparam signed [5:0] p17 = {4{{4{(-2'sd1)}}}};

  assign y0 = ((($unsigned((a1&&a4))&{3{p8}})&&{4{(-b2)}}));
  assign y1 = {{p15,p14,a5},({b5,b1}!=={a3,b4,a4})};
  assign y2 = ((((p4)?(p14>=p4):{p13,p14}))?(-5'sd2):{2{{p15,p5}}});
  assign y3 = $unsigned($unsigned($unsigned($unsigned(($unsigned($signed(((~&p1)&(p11<p7))))>{$unsigned((4'd2)),(p12>>>a4)})))));
  assign y4 = (~&(!((~|(-(~&(!(p17?p15:p2)))))?(~^(+(p8?p15:p13))):(~^(^(a0?p16:p16))))));
  assign y5 = (|{1{{3{({2{p2}}>>(p14>>p15))}}}});
  assign y6 = (|(~&$signed({(((3'd1))?(~|({p14,p6}+(p8<<p10))):(!(&(~&(a3?p10:p16)))))})));
  assign y7 = {$signed({b3,a1}),$unsigned((b0))};
  assign y8 = ((b5?a1:a1)?(-5'sd6):(b4*a0));
  assign y9 = {2{(((a2==a3)===(~a4))|(!(+(5'd2 * b2))))}};
  assign y10 = (((~|(4'sd0))&&({a0,a3,b2}^~{b5,a2,b0}))!==$signed((4'sd7)));
  assign y11 = (|(&(5'sd2)));
  assign y12 = $signed((&(+(+(~p6)))));
  assign y13 = (((a2?p15:p0)<=(~^(p4*p8)))>>>((6'd2 * p1)^~(p4||p11)));
  assign y14 = $unsigned({4{a0}});
  assign y15 = (~&(4'sd4));
  assign y16 = (~^(3'd0));
  assign y17 = (~&(((~^(3'd6)))!==((4'd5)-(-3'sd1))));
endmodule
