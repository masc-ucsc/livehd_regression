module expression_00891(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((-4'sd5)+(3'd1)),(2'sd0)};
  localparam [4:0] p1 = ((~&(-3'sd0))?((-2'sd1)?(2'd2):(3'sd2)):((4'd0)?(-5'sd12):(-2'sd1)));
  localparam [5:0] p2 = (+{(5'sd0),{(-2'sd1)},(^(4'd8))});
  localparam signed [3:0] p3 = (+(~((-5'sd12)==(2'd2))));
  localparam signed [4:0] p4 = (4'sd2);
  localparam signed [5:0] p5 = ((-3'sd1)?(3'd6):(4'd1));
  localparam [3:0] p6 = {4{((2'd3)^(5'd27))}};
  localparam [4:0] p7 = (&{4{(2'sd0)}});
  localparam [5:0] p8 = (&(|(^(&(&((3'sd0)>>(-4'sd4)))))));
  localparam signed [3:0] p9 = {1{{1{((-5'sd13)?(2'd2):(4'sd3))}}}};
  localparam signed [4:0] p10 = {(!(&(~^(&{{(4'sd6),(-5'sd6)},(~^(4'sd1)),(+(-4'sd5))}))))};
  localparam signed [5:0] p11 = (5'd2 * ((3'd4)>>(2'd3)));
  localparam [3:0] p12 = ((((-2'sd1)>(2'd1))?{3{(-4'sd3)}}:{2{(4'sd4)}})+{4{{1{(-3'sd1)}}}});
  localparam [4:0] p13 = (((4'd11)>>(-3'sd2))==((3'd3)?(3'd3):(-2'sd0)));
  localparam [5:0] p14 = (^(!(-((2'd3)-(-4'sd2)))));
  localparam signed [3:0] p15 = ((!(-5'sd15))?(((5'd24)&&(3'sd0))||(-(5'sd4))):(((5'sd9)^(3'd4))==((4'sd7)+(2'd2))));
  localparam signed [4:0] p16 = ((|(2'd0))?(^(-4'sd7)):{4{(-2'sd1)}});
  localparam signed [5:0] p17 = ((~^{(3'd7)})>>>((2'd1)>=(2'd2)));

  assign y0 = {(^(-4'sd0)),{(~^a5)}};
  assign y1 = (((~|b4)+(b0-p1))+(-(p15%a4)));
  assign y2 = (~&(~&((p3-a2)^~{(-4'sd1)})));
  assign y3 = (+((+(&{(|(~|(!a3)))}))?((a5&a4)^{(a1<b3)}):((b1^b3)>>(a2?p13:b3))));
  assign y4 = {1{(({4{p3}}!=(p3>>b0))>$unsigned({2{(a4-b0)}}))}};
  assign y5 = (-{2{(+(p12>=p16))}});
  assign y6 = ((((a2?p16:b0)-(b5)))+((a0>a3)?(b2?b5:a1):$signed(b4)));
  assign y7 = {{(~b5),{3{p1}},{2{p15}}},{(~&p15),(!p10),(~a5)},{{1{a0}},(~|a0),{b3,p13}}};
  assign y8 = ((a4&b1)>$unsigned(a5));
  assign y9 = (((a0^b1)!==$unsigned(a4))>>>((a3<<p14)^~(a0?p11:a4)));
  assign y10 = ({4{b3}}?(a3?p3:a2):(p14|p12));
  assign y11 = (^(({2{(p10>>>p2)}}&((p2^p12)||(|p0)))>>{3{(b4>>>p12)}}));
  assign y12 = (((3'd6)>>(b2?b0:b5))<((5'sd5)^~(a0|b4)));
  assign y13 = (({4{b5}}^{p6,p12,a3})||{{4{p6}},{p15,a3},(b0===b1)});
  assign y14 = (!((|p11)<=(p2||p11)));
  assign y15 = (({(~^a4),$signed(a5),{a3}})?(-3'sd3):(&$signed((~{$signed($signed(b0))}))));
  assign y16 = (~|b2);
  assign y17 = (~&(|(($signed({1{b5}})|(b0>a3))<<(!{3{$unsigned(b0)}}))));
endmodule
