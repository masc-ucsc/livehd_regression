module expression_00266(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd7);
  localparam [4:0] p1 = (({(2'd3),(-4'sd6),(4'sd5)}|(4'sd1))=={((5'd24)^(-2'sd0))});
  localparam [5:0] p2 = {{2{{3{(-2'sd0)}}}},{1{{{(2'd3),(3'd3),(5'sd8)},((-4'sd1)||(4'd5))}}},{{2{(-5'sd11)}},{(-2'sd1),(3'd0),(-3'sd2)}}};
  localparam signed [3:0] p3 = ((5'sd15)<<<(2'd0));
  localparam signed [4:0] p4 = ((^(5'd8))<<<((2'd3)?(5'd14):(3'd1)));
  localparam signed [5:0] p5 = (+(((5'd21)<=(3'sd2))>=((2'sd0)!=(-5'sd0))));
  localparam [3:0] p6 = ((~|(2'd0))?(~&(-2'sd1)):{(2'sd0)});
  localparam [4:0] p7 = ((((-2'sd1)>=(-5'sd15))?((-3'sd3)|(4'sd3)):((5'd16)?(5'd24):(4'd14)))?(((2'd1)>=(-4'sd0))?(6'd2 * (4'd5)):((2'sd0)/(5'sd0))):((~|(5'd30))+(4'd14)));
  localparam [5:0] p8 = {4{{2{(-4'sd4)}}}};
  localparam signed [3:0] p9 = ((~((4'd10)&(2'd0)))==(+(~^(~&(4'sd1)))));
  localparam signed [4:0] p10 = (~(&((^(^(+(~^(~^(4'sd3))))))===((~^(+(-4'sd2)))!==(~^((2'd3)<<(4'sd1)))))));
  localparam signed [5:0] p11 = (^({3{(4'sd2)}}?((5'd31)?(2'd1):(5'd10)):(~^((3'd2)&&(4'sd3)))));
  localparam [3:0] p12 = {{3{{(4'd2 * ((3'd2)+(2'd2)))}}}};
  localparam [4:0] p13 = (&(~|(((~^(-4'sd1))<(|(2'd1)))==(((5'sd5)>>(-2'sd1))===((4'd1)^~(5'd13))))));
  localparam [5:0] p14 = ((|(4'd4))==={(-2'sd0),(-5'sd13)});
  localparam signed [3:0] p15 = {2{{1{(((-3'sd3)?(2'd2):(5'd13))?{2{(4'sd2)}}:(4'd4))}}}};
  localparam signed [4:0] p16 = (-3'sd3);
  localparam signed [5:0] p17 = ((((3'd6)?(-4'sd5):(4'd12))?((5'sd14)&(2'd3)):(~&(-3'sd1)))?(((3'd0)>>(-3'sd2))?(~&(5'd13)):(|(5'd14))):(2'd0));

  assign y0 = {3{(4'd2 * $unsigned((p0<p4)))}};
  assign y1 = (((a3&&a3)+(5'd16))&&{4{p1}});
  assign y2 = (a4<b1);
  assign y3 = (2'sd1);
  assign y4 = (((a2^a5)<<<$unsigned($signed(b5)))===$signed((($signed(b3)==(a3<<b5)))));
  assign y5 = (&(~|(+(2'd3))));
  assign y6 = (4'sd0);
  assign y7 = (5'd2 * (p8>>>p7));
  assign y8 = (|(-(~^a3)));
  assign y9 = (|(((+b1)!==(b5>>>a4))-(&(p10>p9))));
  assign y10 = (5'sd6);
  assign y11 = (-{(~(~&{(2'sd1),(4'd7)})),(3'sd3),{2{(~(3'd0))}}});
  assign y12 = (((+(p11<=b0))<<<((b0&p5)>=(p10>p11)))&((~(~&(b5)))==($signed(a4)===(!a4))));
  assign y13 = {3{((b3>>p15)>=(a0==a1))}};
  assign y14 = ((5'd21)^~(((b1!=a5)===(5'd30))));
  assign y15 = (&(p13));
  assign y16 = $unsigned((~(p3)));
  assign y17 = (!(4'd11));
endmodule
