module expression_00909(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(3'd1),(3'd6),(2'd0)}^~(((4'sd1)?(3'sd3):(-2'sd1))-{(-2'sd1),(5'd12),(3'd7)}));
  localparam [4:0] p1 = (((+(-3'sd0))&{2{(-5'sd2)}})<<(-((+(2'sd1))<=(^(5'd12)))));
  localparam [5:0] p2 = (-3'sd3);
  localparam signed [3:0] p3 = ({(~|(4'd7)),{(5'd10),(3'd7),(5'd31)}}<<<{(|((5'd5)&(-5'sd9)))});
  localparam signed [4:0] p4 = (4'd2 * ((5'd29)!==(5'd20)));
  localparam signed [5:0] p5 = ((5'd13)<<<(-4'sd5));
  localparam [3:0] p6 = (-3'sd1);
  localparam [4:0] p7 = ((^(-((3'd0)?(5'd7):(4'd13))))==(((5'd21)>>>(3'd2))|(^(5'd31))));
  localparam [5:0] p8 = {(3'd6),(-4'sd4),(5'sd3)};
  localparam signed [3:0] p9 = (5'sd2);
  localparam signed [4:0] p10 = (-(~^(~{(2'd2)})));
  localparam signed [5:0] p11 = {4{(-5'sd0)}};
  localparam [3:0] p12 = (((((4'd7)%(4'd7))*((-2'sd1)*(2'd2)))&(((4'sd0)===(5'sd4))!==((2'd1)!=(3'd5))))^((((5'd6)>(-5'sd3))!=((-2'sd1)|(-5'sd6)))<(((4'sd6)<(4'd10))==((3'd5)>>>(5'sd10)))));
  localparam [4:0] p13 = {(~(((2'sd0)>=(2'd0))==((3'd7)>(5'd12)))),{((-5'sd14)>>>(3'sd1)),((4'sd3)>=(5'sd9))}};
  localparam [5:0] p14 = {1{(-(((2'sd0)==(2'd3))!=((4'sd7)>>(4'd15))))}};
  localparam signed [3:0] p15 = (+((-5'sd0)?(~(5'sd10)):((4'd8)<=(-5'sd6))));
  localparam signed [4:0] p16 = (!((((5'sd10)?(4'd0):(3'd5))?(~^(-5'sd13)):(~&(4'd10)))?(&((4'd9)?(2'd3):(5'd27))):((~&(3'sd0))?((2'd0)?(-5'sd15):(-2'sd1)):((2'sd1)?(4'd15):(2'd0)))));
  localparam signed [5:0] p17 = (((6'd2 * (5'd13))<<(~(4'sd2)))<=(|((2'sd0)^~(5'd24))));

  assign y0 = (|(~{(+(|(~{{{(!(~^{a5,a5})),(|(~&(+b5)))}}})))}));
  assign y1 = {(~&(3'd7))};
  assign y2 = (|(~|(-(((~^(p8!=p3))==(|(|{1{p1}})))|(~|$unsigned({3{(5'd2 * p2)}}))))));
  assign y3 = (6'd2 * (p6^b1));
  assign y4 = (($signed((p16<<p2))<=($signed(p0)==$signed(a4)))!=((-4'sd5)>=(3'd7)));
  assign y5 = (+(^(~(!((~^$unsigned((~|(b4))))===((-a0)>>(|a4)))))));
  assign y6 = $signed((^(4'd13)));
  assign y7 = ((3'sd1)>(5'd18));
  assign y8 = (((b3!=p13)?(b5>>a1):(a0>>a4))?((-3'sd3)!==(-4'sd0)):((b1?b0:a5)?(a0!==a3):(4'sd2)));
  assign y9 = ((2'd3)>>{2{$signed(a3)}});
  assign y10 = (~&(((a2!=b3)!==(5'sd12))?(4'sd7):(4'd5)));
  assign y11 = (a1>>>a5);
  assign y12 = {1{({4{p6}}+{2{p11}})}};
  assign y13 = {{{(5'd6),{(a0||a1),{a4,a0}}}},{$signed({(4'd3)})}};
  assign y14 = (({3{p3}}<=(a0===b5))!={1{($signed(b5))}});
  assign y15 = ((p6&&p0)<<<{1{p3}});
  assign y16 = ({p16,p1,a4}>=(-3'sd3));
  assign y17 = {{{b0},{b1,b2,a4},$unsigned(a0)},{{{a3,b5}},$signed($signed(a2))},$signed({{b1},{p10,b0},{b1,a3,a5}})};
endmodule
