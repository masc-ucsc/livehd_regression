module expression_00356(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'sd1)!=(2'd3));
  localparam [4:0] p1 = (~(2'sd0));
  localparam [5:0] p2 = {{(((-3'sd1)==(5'd4))>=((3'd1)||(4'd4)))},({(4'd5)}&&((5'd10)<(4'sd5)))};
  localparam signed [3:0] p3 = ({(4'd3),(2'd1),(2'd1)}<=({(3'd5),(4'sd3),(3'd3)}<<{(2'sd0)}));
  localparam signed [4:0] p4 = ((((4'd11)||(-5'sd10))|{1{((4'd6)!==(5'd7))}})!=={1{(((2'sd0)>=(-4'sd4))+((3'sd1)===(2'sd0)))}});
  localparam signed [5:0] p5 = (((5'sd8)?(2'd2):(-4'sd3))?(&(4'd5)):((2'd0)?(-5'sd10):(5'd6)));
  localparam [3:0] p6 = ((5'd15)<<((5'd19)>>>(|(4'd15))));
  localparam [4:0] p7 = ((-(((3'd5)?(3'd3):(4'd0))>>{(2'd0),(-2'sd0)}))<<(|({(2'd3),(3'd2)}<<(~|(2'd0)))));
  localparam [5:0] p8 = {({(5'd28),(-2'sd1),(3'd2)}^~(&(3'd0))),(6'd2 * (2'd2)),(((2'd2)<(4'd14))-((5'sd1)+(5'd29)))};
  localparam signed [3:0] p9 = (!(-2'sd0));
  localparam signed [4:0] p10 = (^(((&((4'sd2)!==(-5'sd0)))^((3'd5)===(5'd23)))<<(((5'd9)&(4'sd6))>((-4'sd0)>>(5'sd7)))));
  localparam signed [5:0] p11 = ({4{(4'd4)}}^(((-3'sd3)<<<(-3'sd3))<<((3'd0)&(2'sd1))));
  localparam [3:0] p12 = (((2'd0)?(-5'sd9):(-3'sd2))*((3'd3)?(4'd2):(3'd4)));
  localparam [4:0] p13 = (({1{((3'sd0)>>>(-2'sd0))}}==={1{((-5'sd1)^~(3'd4))}})>=(4'd2 * ((3'd3)&(4'd7))));
  localparam [5:0] p14 = {1{(~|{1{{2{(|(4'sd5))}}}})}};
  localparam signed [3:0] p15 = {{3{(3'd3)}}};
  localparam signed [4:0] p16 = ({(4'sd3)}-{4{(4'sd5)}});
  localparam signed [5:0] p17 = ((((3'sd2)>>(-2'sd0))<=(6'd2 * (2'd1)))|(((2'd3)>=(-5'sd13))>((-2'sd1)^(3'd4))));

  assign y0 = {4{b2}};
  assign y1 = (((p13&&p11)>(p4?a3:p0))<=((b1===b4)?(p6%a5):$signed(a5)));
  assign y2 = {(~|{2{{p3,p13}}}),(&{3{(5'd2 * p0)}})};
  assign y3 = ((~^(~|$signed((3'sd0))))<<<((&a3)?(~p13):(^p7)));
  assign y4 = (((p7?a2:b1)?{p15,p1}:{b5})?$unsigned({4{p15}}):$unsigned({(4'd0),(&a0)}));
  assign y5 = {(^(~&((p0<=p11)?{4{p7}}:(b5+p14)))),(!(|((~&(p13<p10))&&(p9^p16))))};
  assign y6 = {4{p16}};
  assign y7 = ($unsigned((^$unsigned($signed((-$unsigned((!b5))))))));
  assign y8 = {({3{a4}}>={1{a1}}),{2{{a0,a3}}},((4'sd7)<<{b0,a5})};
  assign y9 = (({1{{4{(p3)}}}}-$signed({1{{2{(p1-a1)}}}})));
  assign y10 = {{b4,p10},(6'd2 * a0)};
  assign y11 = ((^{(b2!==a0),(b5!==b2),(b3&&a4)})<=$signed({$signed((b2>>>a2)),{(b5>a2)},(~|(+b4))}));
  assign y12 = (($unsigned(p0)?$signed(b3):(p13?p12:b5))>((b5||p1)?(b5):$signed(a2)));
  assign y13 = {(4'sd3),((5'd12)=={1{a5}})};
  assign y14 = {{4{{1{p4}}}}};
  assign y15 = (((p1||p8)+$signed(b4))>({p5,p15}<<(3'd0)));
  assign y16 = ({4{{p9}}}>>((~&{4{p8}})-{p4,p1,p14}));
  assign y17 = ({(p4&p16),(3'sd1),(p3<<p14)}>>((3'd6)^{b5,a0}));
endmodule
