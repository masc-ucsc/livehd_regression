module expression_00024(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(3'd4));
  localparam [4:0] p1 = (((-2'sd1)<<<(3'd3))>((2'd0)<(3'sd1)));
  localparam [5:0] p2 = ({(-3'sd2)}?((5'd22)<<(4'd6)):((5'sd5)>=(2'sd1)));
  localparam signed [3:0] p3 = (~&(2'd2));
  localparam signed [4:0] p4 = ((((2'd1)|(3'sd0))<<<(~|(5'sd4)))>=({(4'sd3),(2'd2),(3'd7)}+(~(3'd1))));
  localparam signed [5:0] p5 = (4'd6);
  localparam [3:0] p6 = ((-3'sd3)?(-5'sd9):(4'd15));
  localparam [4:0] p7 = ((((4'd15)>=(4'd12))&&{(2'd1),(3'd4)})?({(4'd9)}&((4'd4)?(5'sd13):(-3'sd3))):((3'sd3)?(3'd7):((5'd20)^(5'sd15))));
  localparam [5:0] p8 = ((3'sd2)^~(((2'sd0)?(3'd3):(5'sd5))!=((3'sd2)!==(4'd4))));
  localparam signed [3:0] p9 = ({2{{4{(5'sd3)}}}}==((&(4'sd2))?(~|(5'd10)):((3'd1)&(4'd2))));
  localparam signed [4:0] p10 = (&({(5'd19)}?((2'd1)<<<(2'd0)):((4'd6)?(-3'sd0):(-4'sd3))));
  localparam signed [5:0] p11 = (+(^(-(~^(-5'sd7)))));
  localparam [3:0] p12 = (~^(+(~|(5'd5))));
  localparam [4:0] p13 = ((2'sd0)^~(5'sd14));
  localparam [5:0] p14 = (4'sd4);
  localparam signed [3:0] p15 = {(4'd2),((-4'sd1)?(3'sd2):(5'sd5)),(!(3'sd0))};
  localparam signed [4:0] p16 = (~|{1{(~^((5'd31)?(-3'sd2):(3'd3)))}});
  localparam signed [5:0] p17 = (&{{(2'd0)}});

  assign y0 = $signed((5'sd5));
  assign y1 = (-($signed(((~^p10)>>>(p2<p12)))?($signed((p13?p17:p14))>>>(p5?p14:p17)):((p9?p7:p13)+(p6&&p6))));
  assign y2 = {4{{1{{2{p11}}}}}};
  assign y3 = (5'sd8);
  assign y4 = (^((^{1{(p5||p12)}})));
  assign y5 = {4{(3'd4)}};
  assign y6 = (&(-((a1?b1:b1)&(!b3))));
  assign y7 = (((!{$unsigned(p14),(3'sd2)})<=((p3<<<p11)||(4'sd2)))^~(2'd0));
  assign y8 = (^(2'd1));
  assign y9 = (p2<<p4);
  assign y10 = (((a4&&a2)!==(b5?a4:b5))?((b3!=a5)<<(a4!==b4)):{b5,b5,a1});
  assign y11 = ((b3<b0)<(a2&p12));
  assign y12 = ({4{b3}}^~$signed((a0<b2)));
  assign y13 = (&($signed((^$unsigned(((2'sd1)!=(b2<<b2)))))!==((~&($signed((2'd0))>>$signed((~a5)))))));
  assign y14 = (-5'sd7);
  assign y15 = {(!{(2'd1),(~&{b3,p4})})};
  assign y16 = ($signed((3'sd3)));
  assign y17 = ((((p16/b1)<<(a0<<<p13))^((a3||p6)+(p8<<<p15)))|(((p0<p15)>>>(4'd2 * p7))||((p13-p14)&(b1^p9))));
endmodule
