module expression_00442(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd0);
  localparam [4:0] p1 = (~&(~|(~&(-(~|({(3'd1),(2'sd0),(5'd19)}^((3'sd1)||(5'd31))))))));
  localparam [5:0] p2 = (-2'sd1);
  localparam signed [3:0] p3 = (&(~^(&(2'd3))));
  localparam signed [4:0] p4 = (5'd13);
  localparam signed [5:0] p5 = ({4{(2'd2)}}!=({1{(5'd21)}}+((2'sd0)?(2'd0):(5'sd9))));
  localparam [3:0] p6 = ((-(4'd12))+(-2'sd0));
  localparam [4:0] p7 = {2{((-2'sd1)<<(3'd5))}};
  localparam [5:0] p8 = {1{((2'd2)>=(-4'sd7))}};
  localparam signed [3:0] p9 = {{(4'd11),(-4'sd6)},((2'sd1)&(4'sd7)),((4'd10)?(2'sd0):(3'd5))};
  localparam signed [4:0] p10 = ((-2'sd0)?(3'd7):(3'd5));
  localparam signed [5:0] p11 = ((((-2'sd0)%(2'd3))||((4'sd5)|(2'sd1)))||(((5'd29)+(5'd31))!=((4'sd1)?(-4'sd6):(3'd7))));
  localparam [3:0] p12 = ({2{(-4'sd5)}}<<<(+{1{(~(!((3'sd2)>(5'sd12))))}}));
  localparam [4:0] p13 = (|(~(~&(~&(-(&(~(-(&(&(~&(!(3'sd2)))))))))))));
  localparam [5:0] p14 = ({4{(3'd6)}}==(^(5'sd10)));
  localparam signed [3:0] p15 = ({2{{3{(-2'sd1)}}}}!==({2{(5'd6)}}<<((2'sd1)>=(4'd9))));
  localparam signed [4:0] p16 = ({4{(2'sd1)}}||(4'd13));
  localparam signed [5:0] p17 = (~&(-4'sd3));

  assign y0 = (($unsigned((b3===a5))>{$signed(b3)})-((b4)?(b1):(2'd3)));
  assign y1 = (!({3{(&$signed(p0))}}>(-{4{(p15)}})));
  assign y2 = {4{(~|(b0<<<b4))}};
  assign y3 = (((p11^a0)<=(4'd3)));
  assign y4 = (!(4'd0));
  assign y5 = (3'd3);
  assign y6 = {1{(!((~|{1{a0}})?(b3==p12):(^{p16,b1,b2})))}};
  assign y7 = (~|(+(|(((a1!==b4)===(b2>=b4))>>((p15>=p13)|(~&(~^p0)))))));
  assign y8 = $signed((&(~|(~&((~p12)?(a0):(a5<b1))))));
  assign y9 = (((a5^~a0))===$unsigned(((a3<<b2))));
  assign y10 = {({3{b5}}<=(&(~^{2{p17}})))};
  assign y11 = ({a0}<(b5?a5:b2));
  assign y12 = (2'd0);
  assign y13 = (2'sd0);
  assign y14 = ({3{(b1||b2)}}>(5'd2 * (5'd1)));
  assign y15 = (!(-5'sd8));
  assign y16 = (3'd6);
  assign y17 = (~&(((~^(~&(~|p17)))>>>((a2!==a5)!=(b4<p1)))<(((b0!==b0)+(!p5))+(!(~(~^p2))))));
endmodule
