module expression_00910(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd7)||((5'd6)<<(4'd2)));
  localparam [4:0] p1 = (4'd8);
  localparam [5:0] p2 = (~^((2'd0)<{1{(&(5'd25))}}));
  localparam signed [3:0] p3 = ((2'd3)?(4'd6):(-5'sd2));
  localparam signed [4:0] p4 = {2{(-2'sd0)}};
  localparam signed [5:0] p5 = (-3'sd3);
  localparam [3:0] p6 = ((((5'sd4)<<(3'd2))>(3'sd3))>>>(-(-(!(3'sd0)))));
  localparam [4:0] p7 = (+(~&(!(|((3'd3)<(4'd7))))));
  localparam [5:0] p8 = ((^((-5'sd13)!==(2'd1)))^~((-(5'sd15))===((4'd8)?(3'sd0):(5'd3))));
  localparam signed [3:0] p9 = {(-(2'sd0)),((3'd7)===(4'd12)),(2'd2)};
  localparam signed [4:0] p10 = (~&(~^(&(~&(^(+(~^(!(~(+(~^(~(!(~(5'd5)))))))))))))));
  localparam signed [5:0] p11 = ((~|{(+(!(2'sd1))),((5'd18)?(5'd1):(-2'sd0))})<<<(((-3'sd0)?(5'd26):(4'd5))?((4'd11)?(-4'sd0):(4'sd0)):{1{{4{(4'sd7)}}}}));
  localparam [3:0] p12 = ((3'd3)?(4'd1):(5'd24));
  localparam [4:0] p13 = (((2'sd1)?(3'sd3):(-5'sd12))!=((5'd25)^(-5'sd6)));
  localparam [5:0] p14 = {{{(4'sd1),(4'd5)},(((2'd0)>>(2'sd0))>>>((2'd2)<<(4'd14)))}};
  localparam signed [3:0] p15 = (((4'sd7)?(-2'sd1):(3'd5))?((-5'sd15)<(2'sd1)):((3'd2)&(-2'sd1)));
  localparam signed [4:0] p16 = (~((|(~|((!(5'sd7))==(~&(-2'sd0)))))^~(~&(|(+((4'd14)&(5'sd1)))))));
  localparam signed [5:0] p17 = (2'd3);

  assign y0 = (3'd6);
  assign y1 = (((a2?b4:a3)?(b3|a1):(b1<<b0))===($signed(b3)?(-a4):(a2?a5:b4)));
  assign y2 = (3'd0);
  assign y3 = (~&{4{p0}});
  assign y4 = {($unsigned({2{p15}})^{p17,p5,p5}),$signed(({1{a5}}!==$unsigned(b3)))};
  assign y5 = (((~&((p1+p10)!=(p13^p17)))>>>((p7/p0)!=(p4%p3)))<=(((p17>>>p5)<=(|p3))>=((!p2)+(&p11))));
  assign y6 = (((3'd5)-(p9|p3))?(4'd2 * (p6<p7)):(4'd3));
  assign y7 = (((p10?p13:p3))==(p6>>>p2));
  assign y8 = ((~((~(a1>>b5))>>{b4,b2}))!==(6'd2 * (-(b1>>>b1))));
  assign y9 = (~(-{(2'sd0),(p1>>>b2),$signed(b3)}));
  assign y10 = (5'd20);
  assign y11 = (!(&(~|(3'd6))));
  assign y12 = ({({{b1,a5,b0},(b5===a5)}<<<((b2<<<a2)===(a3>>>a1)))}^~{({(b0!=a2),{a5,a5}}+({b0}&&(a5!==b2)))});
  assign y13 = (-{3{(-2'sd0)}});
  assign y14 = ({(a3!==a4),(b0?b1:p9)}?((4'd2 * p2)?{b3}:(b3?a5:a0)):{{a2},(a2?a1:a5),{b5,a5}});
  assign y15 = (&(&$signed((a3?a1:a2))));
  assign y16 = (~^(-((!{(p4>=p12),{p2,p12,p10},(!p9)})&((p16^~p7)<<<(|(p16==p16))))));
  assign y17 = ((~^(+a1))!=(p2*p3));
endmodule
