module expression_00696(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(-2'sd0)}};
  localparam [4:0] p1 = (({1{(5'sd7)}}^~((2'd0)!=(2'd3)))<((2'd2)>>>((3'd4)!==(4'd4))));
  localparam [5:0] p2 = ((((5'd14)^(2'sd1))?((4'd6)*(-5'sd15)):((-2'sd1)<=(3'sd2)))|((|(4'd13))|(2'd0)));
  localparam signed [3:0] p3 = (5'sd3);
  localparam signed [4:0] p4 = ((2'sd0)===(-2'sd1));
  localparam signed [5:0] p5 = (((~|(-4'sd3))<(-(3'sd3)))-(5'd2 * (~&((2'd0)|(4'd15)))));
  localparam [3:0] p6 = (&(-(-(((2'sd1)?(2'd3):(3'd3))?((3'd1)?(5'd8):(5'd14)):((2'd2)?(2'sd1):(-4'sd6))))));
  localparam [4:0] p7 = {((4'sd0)>(2'd3)),((3'sd0)?(2'd2):(4'd6))};
  localparam [5:0] p8 = (~(3'sd2));
  localparam signed [3:0] p9 = {4{{4{(3'd0)}}}};
  localparam signed [4:0] p10 = (~(2'd2));
  localparam signed [5:0] p11 = (~|(~^((5'sd13)?(-3'sd3):(-4'sd2))));
  localparam [3:0] p12 = ((((-2'sd0)&(2'sd0))+((2'sd0)&(-5'sd10)))&(2'd1));
  localparam [4:0] p13 = (-(3'd7));
  localparam [5:0] p14 = ((5'sd4)?(-5'sd8):(-3'sd2));
  localparam signed [3:0] p15 = ((|(5'd30))||{(2'sd0),(2'd0)});
  localparam signed [4:0] p16 = (~(~((-((5'sd4)-(4'sd6)))^(~(-(!(-5'sd11)))))));
  localparam signed [5:0] p17 = (!(2'd0));

  assign y0 = ($signed(((((a1>p12)))|((a3^p7)!=$unsigned(p16))))&(((a3>>>p12)&&$unsigned(a1))>=((b4<=p10)<<<$unsigned(p15))));
  assign y1 = ({p12}<=(p12?p14:p3));
  assign y2 = ({(a0-a1),(-b2),(+b4)}!=(-((6'd2 * b0)===(~b5))));
  assign y3 = ((-{{a0,b4},(a1|b4),(b5&a1)})===(~&((^(^a4))&(a0==a2))));
  assign y4 = $unsigned((({p12,p6,p0}&&(~|p5))));
  assign y5 = ((p2|p7)?(p11):(p4?p3:p17));
  assign y6 = (-5'sd15);
  assign y7 = (p6?p1:p7);
  assign y8 = (~&(-3'sd1));
  assign y9 = $signed(($signed(({4{b2}}+(p13!=b1)))));
  assign y10 = $signed((a3?b4:p0));
  assign y11 = ((b4?a0:p8)?(b3?b0:a5):(~p17));
  assign y12 = ({b1,p12,p4}||(4'd2 * (4'd7)));
  assign y13 = (a4?a1:p16);
  assign y14 = ((-4'sd4)?(b2?b2:p0):(-4'sd6));
  assign y15 = (&{(((p3-p2)-$signed(b3))>=({(&a0)})),((+(3'sd3))+(2'd2))});
  assign y16 = (-{3{(&({1{(&(~^p7))}}))}});
  assign y17 = ((3'sd3)?((b0?a0:b2)?{p6,b2,b0}:(-2'sd1)):(3'd5));
endmodule
