module expression_00178(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(((3'sd3)?(-3'sd2):(5'd26))+(|(4'd8))));
  localparam [4:0] p1 = {(~&({(4'sd0),(2'd0)}!=(3'd0))),(~^((~&(3'd5))&(~(5'd16))))};
  localparam [5:0] p2 = ((!(|(2'd1)))*(&((4'd14)*(-5'sd8))));
  localparam signed [3:0] p3 = ((4'd15)>>(2'sd0));
  localparam signed [4:0] p4 = {3{({(-4'sd7),(-2'sd0),(-5'sd4)}<=((5'd5)&(-5'sd11)))}};
  localparam signed [5:0] p5 = (~&(!{2{({1{(4'd5)}}+((2'd0)<=(2'd2)))}}));
  localparam [3:0] p6 = (~(&((+(-4'sd7))?(+(-5'sd14)):((2'sd1)?(5'd9):(3'd3)))));
  localparam [4:0] p7 = ((((-3'sd3)?(3'd1):(2'd2))?(~^(+(4'd13))):((-2'sd1)%(4'sd2)))|(~|(((2'sd0)^(-2'sd1))>((-2'sd0)*(2'd1)))));
  localparam [5:0] p8 = (((2'd1)>=(3'd4))<((2'd3)!=(5'd20)));
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = {{1{(!{{(3'sd0),(3'd5),(5'sd6)},(~&(-3'sd0)),{1{(3'd6)}}})}},(((5'sd4)===(3'd5))|((5'd29)^~(4'd15)))};
  localparam signed [5:0] p11 = (((3'd5)%(5'd25))?(&((-2'sd0)?(3'd3):(4'd5))):(5'd2 * (3'd1)));
  localparam [3:0] p12 = {4{((5'sd8)?(-3'sd0):(3'sd0))}};
  localparam [4:0] p13 = {4{{1{((3'sd3)&(4'sd0))}}}};
  localparam [5:0] p14 = (~&(-5'sd8));
  localparam signed [3:0] p15 = ({4{(-2'sd0)}}-(((3'sd2)>>(4'd10))<=((5'sd6)^(5'd22))));
  localparam signed [4:0] p16 = ((|{1{(!(-5'sd4))}})&&(&(~(^{3{(3'sd3)}}))));
  localparam signed [5:0] p17 = {3{(5'sd9)}};

  assign y0 = {(-(5'sd12)),(3'sd0)};
  assign y1 = (((2'sd1)==((-4'sd7)!=(|p15)))>>>(~&(~|((b0^~b2)<<<(-4'sd6)))));
  assign y2 = ((b1/p2)<=(-5'sd3));
  assign y3 = {{3{p10}},(4'sd4),({a5,a3,b5}==={1{a2}})};
  assign y4 = {2{(|(~|(-2'sd1)))}};
  assign y5 = (a3>>>a0);
  assign y6 = {((a5&a1)^(!{2{a3}})),{1{{3{(b1?b5:b5)}}}},({a0,p0,b3}?{2{b0}}:{b1,b4})};
  assign y7 = (((b1>a1)?$signed(a5):(b2>>a2))^~(-((5'd2 * a2)-$signed(a3))));
  assign y8 = {1{(((-3'sd3)===((4'sd1)<<(b2<a4)))!=(((-2'sd0)<=(a0>a5))|((a0^~b3)-{3{b0}})))}};
  assign y9 = {3{(p11?p14:p16)}};
  assign y10 = (({1{(p10<<<b4)}})+({1{b5}}!==(a4!==a1)));
  assign y11 = {1{(2'd1)}};
  assign y12 = ((4'd6)|(3'd3));
  assign y13 = {2{{(|p13),{3{p1}},{3{p2}}}}};
  assign y14 = {{p5},(&p10)};
  assign y15 = (((p11?b0:a2)!=(|(b5?p0:b1)))-({4{p9}}^(p15?a5:b3)));
  assign y16 = ({2{b5}});
  assign y17 = ({1{((p6?p15:a1)?(p12?p13:p7):{4{a1}})}}|{4{(p10&&b5)}});
endmodule
