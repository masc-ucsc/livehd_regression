module expression_00134(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{{4{(^(4'd3))}}}};
  localparam [4:0] p1 = ({1{{2{(5'd27)}}}}-({4{(2'd0)}}|((3'd0)||(-5'sd6))));
  localparam [5:0] p2 = {{(4'd2),{(2'd2),(4'sd4),(-5'sd10)}},(^(+(2'sd1))),(3'sd1)};
  localparam signed [3:0] p3 = (5'd19);
  localparam signed [4:0] p4 = (((3'sd2)!==(5'sd8))*(|(~&(3'sd2))));
  localparam signed [5:0] p5 = {({(5'd29),(3'sd0)}==={(2'd0),(3'sd3),(3'd0)}),(((3'sd2)||(5'd26))-{(4'd5),(2'd3)})};
  localparam [3:0] p6 = (&(2'd3));
  localparam [4:0] p7 = (~|(((4'sd7)%(5'd4))*(~^(5'd30))));
  localparam [5:0] p8 = (^(5'sd5));
  localparam signed [3:0] p9 = {3{((5'sd0)>>(3'sd1))}};
  localparam signed [4:0] p10 = (((3'd3)?(-4'sd2):(2'd3))?((-(4'sd5))&&((5'd31)!=(3'sd2))):(((3'd3)>>(3'd2))<((-3'sd0)&&(2'd2))));
  localparam signed [5:0] p11 = ((-3'sd0)&&(5'd2 * (5'd12)));
  localparam [3:0] p12 = {(~&(&(-3'sd3))),(+(|(-3'sd1))),(|(^(5'd20)))};
  localparam [4:0] p13 = (~|(2'sd1));
  localparam [5:0] p14 = {({{(5'sd9),(4'd0)},((5'd0)<=(-2'sd0))}&(-{(+(4'sd0))}))};
  localparam signed [3:0] p15 = ((5'd2 * ((2'd2)*(3'd7)))===(((-5'sd10)<<<(3'd0))^((4'd3)|(3'd7))));
  localparam signed [4:0] p16 = (((-2'sd1)?(2'd0):(3'sd2))?{2{{(5'd30)}}}:({1{(2'd2)}}<=(-4'sd5)));
  localparam signed [5:0] p17 = (2'd3);

  assign y0 = $unsigned($signed(($unsigned($unsigned(($signed(($unsigned($unsigned(($unsigned($unsigned($unsigned($signed(p14)))))))))))))));
  assign y1 = $unsigned(((~^(p9==p2))&&(^(p12?p6:p4))));
  assign y2 = ({((p12-p12)<<{2{p8}})}<((p7>=p7)-$unsigned((a3==p3))));
  assign y3 = (((b2?b2:b1)&&(b5?p9:a5))>((a2===a0)==(^{2{a2}})));
  assign y4 = ($unsigned((b4===a3))!=(4'd2 * b1));
  assign y5 = {((|b2)?(p2?a1:b1):(a5<b2)),{(-3'sd3),(~|b2),(3'sd3)},(&{(4'd10),(a4>>b5)})};
  assign y6 = (((b3<<<p6)^(b5&a0))&((b0>>>a5)&&$signed({a3,a1,p15})));
  assign y7 = (((p9!=b2)>>{1{(5'd25)}})>>>({3{b3}}>=(~(b0<=b3))));
  assign y8 = ($signed(((4'd3)))?$signed(((4'd4)?(4'd4):$unsigned(b0))):(3'sd3));
  assign y9 = ({4{(~&a4)}}?((~^(b4<<a3))&(~(b4?a3:b0))):((b3>>a2)+$signed((5'd23))));
  assign y10 = ((b5?a3:p12)?(p5?p13:a2):(b3>>p3));
  assign y11 = ((!((~p10)^(p9==p11)))<=(~&(!((~p13)&(~|p15)))));
  assign y12 = {3{$unsigned(((b2>>>p0)))}};
  assign y13 = ($unsigned({1{((a1?b0:a1))}})===(4'sd5));
  assign y14 = (5'd2 * (&(b0+a0)));
  assign y15 = (5'd21);
  assign y16 = (-4'sd0);
  assign y17 = (~^(-5'sd10));
endmodule
