module expression_00105(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|((5'd2 * (!(3'd6)))?(~(5'sd7)):(5'sd8)));
  localparam [4:0] p1 = ((2'd1)!=(-4'sd5));
  localparam [5:0] p2 = ({(-5'sd9)}?((4'd6)?(-2'sd1):(2'd1)):((3'sd3)?(-2'sd0):(3'd3)));
  localparam signed [3:0] p3 = (((4'd0)?(-4'sd7):(5'd26))?(((5'd19)!=(3'd4))>=((5'd26)&(2'd1))):({3{(3'sd1)}}!=={4{(2'd3)}}));
  localparam signed [4:0] p4 = (((-2'sd0)&&(2'd2))?((2'd0)^(3'sd2)):((4'sd3)^(-5'sd3)));
  localparam signed [5:0] p5 = (^((5'd14)?(-2'sd1):(5'd22)));
  localparam [3:0] p6 = {2{{((-5'sd2)&&(5'd16)),((2'd3)|(3'd5))}}};
  localparam [4:0] p7 = {4{{4{(2'sd1)}}}};
  localparam [5:0] p8 = (~(2'd0));
  localparam signed [3:0] p9 = (+(5'd30));
  localparam signed [4:0] p10 = {({3{(5'd25)}}?((-2'sd0)==(3'sd3)):{(3'sd0),(3'd4)}),(3'sd2)};
  localparam signed [5:0] p11 = ((-3'sd0)<<(|((3'sd0)/(5'd13))));
  localparam [3:0] p12 = ((-3'sd1)^~(4'd11));
  localparam [4:0] p13 = ((((3'd0)?(2'd3):(3'd4))?((2'sd0)-(-3'sd1)):((2'd1)<<(-3'sd3)))+(((4'd14)<(-5'sd6))<<((5'd14)>(2'd0))));
  localparam [5:0] p14 = ((((3'sd2)!==(-4'sd0))-((2'd2)?(4'sd0):(4'd13)))>(((-3'sd3)>>(2'sd0))||((-5'sd14)-(4'sd2))));
  localparam signed [3:0] p15 = ((+({3{(-4'sd0)}}&&{(2'd0),(2'd3)}))?(|(~&(|{(2'd2),(3'd5),(5'sd14)}))):(((3'sd3)<(3'd3))>(~^(4'd6))));
  localparam signed [4:0] p16 = (~&(|(6'd2 * ((2'd0)||(3'd4)))));
  localparam signed [5:0] p17 = {2{({4{(-3'sd0)}}||{4{(5'd2)}})}};

  assign y0 = {4{(p16&b5)}};
  assign y1 = ({(b1>a3)}<(~&(b0|a1)));
  assign y2 = (((~|$signed((($unsigned(p14)<(5'd2 * p2))))))^~(((~&p12)||(p14*p14))^$signed((!(^p10)))));
  assign y3 = {3{{1{{2{{3{b4}}}}}}}};
  assign y4 = {2{(((!b0)^(a1>p14))&&((b2?a5:a5)||{2{p16}}))}};
  assign y5 = (2'd1);
  assign y6 = (((p3?b0:p1)?(4'd4):{2{a5}})?({4{p12}}?(b0|p10):(b2?b2:a2)):{1{(2'd0)}});
  assign y7 = $unsigned({$signed({4{p7}}),{(p14+p10),{1{a4}},(b0===a0)},{2{$signed(p17)}}});
  assign y8 = ((^{3{{p1,p13}}})?{(+(p7?p2:p6))}:{4{(|p1)}});
  assign y9 = ({2{{2{b4}}}}||{({1{(b5||p7)}}<=(b0>b2))});
  assign y10 = (5'sd6);
  assign y11 = (3'd5);
  assign y12 = {(+b2),(|p10),(-b5)};
  assign y13 = {2{{1{(5'd2 * (p6!=a1))}}}};
  assign y14 = $signed((a5?p17:p17));
  assign y15 = (p7?p6:p5);
  assign y16 = ((((a4>>p15)<<(3'sd2))^~(-3'sd3))>>(3'sd1));
  assign y17 = ((3'd6)?$signed(p1):{b4,a5});
endmodule
