module expression_00540(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(-{4{((4'd5)?(-3'sd2):(4'd8))}})}};
  localparam [4:0] p1 = (((4'sd0)==(-5'sd6))||{4{(-4'sd3)}});
  localparam [5:0] p2 = (!((2'd3)?(3'sd1):(3'sd3)));
  localparam signed [3:0] p3 = (&(&(-{{(2'sd1),(5'd11)}})));
  localparam signed [4:0] p4 = (&{1{(((-4'sd3)&(-4'sd7))!=(!((3'd4)+(4'sd5))))}});
  localparam signed [5:0] p5 = (4'd5);
  localparam [3:0] p6 = (((3'd3)?(5'd11):(-4'sd7))<=((5'd23)|(5'd5)));
  localparam [4:0] p7 = (((5'd17)?(4'sd3):(5'd27))?((-2'sd1)%(4'd11)):((2'sd0)+(4'sd5)));
  localparam [5:0] p8 = ({(2'sd1)}&((2'd2)>=(4'd12)));
  localparam signed [3:0] p9 = (-3'sd2);
  localparam signed [4:0] p10 = {1{((4'sd3)>=(4'd11))}};
  localparam signed [5:0] p11 = (|{(~&(~|{3{{2{{(3'sd0),(5'd3),(5'd20)}}}}}))});
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = (-3'sd3);
  localparam [5:0] p14 = (~&{(!{((-5'sd12)?(-2'sd0):(-2'sd0)),((5'sd5)&(-5'sd12))})});
  localparam signed [3:0] p15 = (((-4'sd1)?(-2'sd0):(2'sd1))?(-5'sd12):((-4'sd1)?(-5'sd8):(5'sd7)));
  localparam signed [4:0] p16 = {(3'd0),(-4'sd4),(2'd0)};
  localparam signed [5:0] p17 = (-2'sd1);

  assign y0 = {2{(~&($unsigned((b3||b4))&&(b1?b0:p4)))}};
  assign y1 = {1{{(p6<<<p4)}}};
  assign y2 = (a3<<b1);
  assign y3 = ((^a4)?(p1==p9):(|p12));
  assign y4 = {2{(|(~&{2{(~&(|b0))}}))}};
  assign y5 = (({4{p3}}?(-5'sd9):(p12?p12:p9))?((~|p6)?{3{p6}}:(5'd13)):((~p16)&(2'd2)));
  assign y6 = (~^((|(5'sd9))));
  assign y7 = (((p1<<b0)&(p3-p10))!=(2'sd1));
  assign y8 = (3'sd3);
  assign y9 = (~(^(&(~(+(~^(-(-(^(~&(~|(~^(&(^(^p13)))))))))))))));
  assign y10 = (({3{a0}}&&(a0?a0:b2))?((b5<<b0)&&(b2&a3)):{3{(a3>>>a1)}});
  assign y11 = ({(-2'sd0)}!=((4'd11)));
  assign y12 = (p13==b0);
  assign y13 = (+(5'd14));
  assign y14 = ({(&p15),(!p0)}==((p7>>>b0)<(-5'sd0)));
  assign y15 = (({(p17^p16)}<=(p15?p11:p4))>={{p2,p1},{p0,p3,p4}});
  assign y16 = (+(-2'sd1));
  assign y17 = {2{(6'd2 * (p0^p1))}};
endmodule
