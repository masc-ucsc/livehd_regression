module expression_00812(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((5'sd13)||(4'sd7))!=(2'd1))?(5'd2 * {(2'd2),(4'd1),(4'd4)}):((4'd1)<={(-2'sd0),(-4'sd4),(2'd3)}));
  localparam [4:0] p1 = (~|((~((5'd29)?(-3'sd3):(-5'sd7)))^~((-4'sd1)%(-5'sd4))));
  localparam [5:0] p2 = (-(!(~{1{(-(~{1{{4{(5'd1)}}}}))}})));
  localparam signed [3:0] p3 = ((2'd3)!==(2'd1));
  localparam signed [4:0] p4 = (-2'sd0);
  localparam signed [5:0] p5 = (-2'sd0);
  localparam [3:0] p6 = {1{({1{((2'd2)?(5'd10):(5'sd14))}}?(~{(5'd25),(-2'sd0),(-3'sd0)}):(-((-4'sd4)>>>(2'd3))))}};
  localparam [4:0] p7 = ((~&((-4'sd0)?(3'sd2):(-3'sd0)))?((-5'sd9)?(3'd7):(2'd0)):(!((3'd3)?(-5'sd1):(4'd6))));
  localparam [5:0] p8 = (~|(&(-5'sd14)));
  localparam signed [3:0] p9 = (-3'sd2);
  localparam signed [4:0] p10 = (((4'sd7)<<(2'sd0))%(2'd2));
  localparam signed [5:0] p11 = ({4{(!(3'sd1))}}^(^({2{(4'd12)}}?((-4'sd4)?(2'd3):(3'sd3)):(~(4'sd3)))));
  localparam [3:0] p12 = ((^(2'sd1))-(((4'd11)?(5'sd5):(2'd3))>((4'd9)>(4'sd4))));
  localparam [4:0] p13 = (({(-5'sd8),(5'd20),(5'sd6)}+(~&(4'sd5)))=={(-2'sd1),(4'd3),(-5'sd5)});
  localparam [5:0] p14 = (-(!((5'd11)>=(3'd0))));
  localparam signed [3:0] p15 = ((((3'd2)^~(4'd5))&&((4'sd0)<<(3'sd0)))&(((3'd4)<<<(-2'sd1))?((2'sd0)<<<(4'sd3)):((5'd15)>(4'sd4))));
  localparam signed [4:0] p16 = (2'd3);
  localparam signed [5:0] p17 = (-(&(5'sd5)));

  assign y0 = ((p1<<b1)+(b1>>p12));
  assign y1 = (($unsigned({3{b1}})<{2{p14}})<$unsigned((~&$unsigned({p3,b0,p16}))));
  assign y2 = {4{((|p14)<<(-4'sd3))}};
  assign y3 = (((a2^~b2)?{(a1?a4:a1)}:(a1>b3))^~((b4?b0:p16)!={b2,a2,b0}));
  assign y4 = ({1{(6'd2 * (4'd4))}}^~{1{(3'd7)}});
  assign y5 = {{3{(&(~^p0))}}};
  assign y6 = $unsigned((&(((a3))|(b3===a3))));
  assign y7 = (((3'd7)^~($signed((a5&a5))))+(((a4&&b1)|(-4'sd4))>>$signed(((a2)<<$signed(a3)))));
  assign y8 = (((p3&&a4)/a5)+(((b2*b1)<<(b5+b0))^((b3!=p7)!=(6'd2 * b1))));
  assign y9 = $unsigned((((a4*a1)!=(|(a2<<<b0)))===$unsigned(((5'd27)^~(3'd0)))));
  assign y10 = {({b5,b4,p14}+(p15<<<p4))};
  assign y11 = (4'sd0);
  assign y12 = ({3{b5}}^(b1==b0));
  assign y13 = (&{4{(b5&p9)}});
  assign y14 = {3{{2{(4'd2 * p12)}}}};
  assign y15 = (((b5-b4)||(b3===a3))^~((b4&&b0)));
  assign y16 = ((((p0||b5)-(a1))<<(+{3{a1}}))==$signed($signed((~|({3{b0}}<<<(a4>>p13))))));
  assign y17 = (((+((b2<<<a0)===$signed(a0))))?(|$signed({1{(a5?a3:b4)}})):((a4===a2)<=(&(~a5))));
endmodule
