module expression_00826(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd8)?(4'sd2):(3'd4))&&(5'sd5))?(-2'sd1):(((3'd1)*(-2'sd1))&((2'd0)===(-5'sd13))));
  localparam [4:0] p1 = (((|(~(5'sd3)))||(3'd5))<(2'd0));
  localparam [5:0] p2 = (^((~|({(-4'sd4)}==(3'd5)))=={(~{1{(5'd18)}}),{(3'd5),(3'sd1)}}));
  localparam signed [3:0] p3 = (&((5'sd11)!==(+(((-5'sd14)===(-2'sd1))>=(|(~(2'd2)))))));
  localparam signed [4:0] p4 = ((-((2'sd1)^~(-3'sd1)))^~((3'sd0)<<<(-3'sd0)));
  localparam signed [5:0] p5 = (+{((~^(2'd1))!==(~|(4'sd1))),{(^(~|(-(-4'sd4))))},{{{(3'd0),(2'd2)}}}});
  localparam [3:0] p6 = (3'd2);
  localparam [4:0] p7 = {((|(4'd2 * (3'd3)))^~(+{(3'd1),(-5'sd13),(2'd3)}))};
  localparam [5:0] p8 = ((4'd3)^(-4'sd1));
  localparam signed [3:0] p9 = ({(4'd11),(5'd22),(4'd0)}^{(3'sd2)});
  localparam signed [4:0] p10 = ((((3'd4)<<<(-4'sd0))^((5'sd0)!=(3'd2)))!=(((2'd0)|(3'd4))&((4'd15)&(2'sd1))));
  localparam signed [5:0] p11 = {2{{2{{3{(5'd13)}}}}}};
  localparam [3:0] p12 = {{(2'sd1),(3'd5)}};
  localparam [4:0] p13 = ({3{((3'd7)?(4'sd7):(3'd1))}}|{{2{(2'd0)}},{{4{(5'd16)}}}});
  localparam [5:0] p14 = (((-3'sd3)||(3'sd0))?((2'd2)<<(3'd0)):(!(3'd1)));
  localparam signed [3:0] p15 = (-3'sd3);
  localparam signed [4:0] p16 = {3{((6'd2 * (5'd22))>>{2{(-2'sd1)}})}};
  localparam signed [5:0] p17 = (((5'd3)%(5'd25))?(((2'd0)&(-5'sd9))?(3'd7):((5'sd15)&(-5'sd13))):(-((4'd10)&&((3'sd1)!==(2'sd1)))));

  assign y0 = (~(({1{p17}}<(!p6))-(&(p3&p3))));
  assign y1 = (+({{a1,b3,b1},{a0,b2},$unsigned(b1)}===({{(a0>>a5),(b2||b4),(a3>=b1)}})));
  assign y2 = (~&(!(5'd16)));
  assign y3 = (((a3>>>a0)?(5'd2 * a0):(b4?a5:b2))!==((a5?b5:a4)===(a3?a4:a1)));
  assign y4 = (-(2'sd1));
  assign y5 = (4'd2);
  assign y6 = {1{(!(|{4{{2{p11}}}}))}};
  assign y7 = $unsigned((((p1<p1)>>>(a1!==a5))<($unsigned((p2))<<(p13%p9))));
  assign y8 = ((a3?p16:p11)?(b1>>p7):(a2<=p8));
  assign y9 = {(~|($signed((b3!==b5))>{(a2&&p16),(p6>>>a1)})),({1{{1{{4{p3}}}}}}>>>$unsigned((^(~(a2|a1)))))};
  assign y10 = (((2'd3)^~(~&(b1<<<a2)))!==((+(a4<<<b4))|(&(~|(4'sd2)))));
  assign y11 = {{{p13},(-p4),(p10<=p1)},({(p8<p4)}==(~{p10,a0})),(~^{(~&(~&(p4+p15)))})};
  assign y12 = {(~&{1{(~^(-p15))}})};
  assign y13 = (p7?b4:p16);
  assign y14 = (({3{b0}}?(p10^a4):(b3>=b3))|(2'd1));
  assign y15 = (~(^(^b0)));
  assign y16 = (5'd2 * (!$unsigned(p9)));
  assign y17 = (((p13&&b4)*(~|(a5%a4)))!=((b1>>b4)>>>(~^(p8^p6))));
endmodule
