module expression_00670(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|{3{{3{(3'd1)}}}});
  localparam [4:0] p1 = {(((5'd11)>=(2'd2))^~{(5'd31),(2'd1),(-5'sd11)}),{(((5'd14)|(-4'sd0))&((-2'sd1)^(4'd3)))}};
  localparam [5:0] p2 = ({(3'sd3),(4'd12),(3'sd3)}!=(6'd2 * (+(2'd2))));
  localparam signed [3:0] p3 = ((&(-3'sd1))!==((-2'sd1)?(3'd4):(5'sd5)));
  localparam signed [4:0] p4 = (-5'sd1);
  localparam signed [5:0] p5 = {({2{(-5'sd9)}}!=((4'sd7)<(2'd3))),{1{((4'sd4)+(2'sd0))}}};
  localparam [3:0] p6 = ((-4'sd2)|(3'd4));
  localparam [4:0] p7 = (+(((-2'sd0)|(-2'sd1))&((2'd1)<<<(4'd0))));
  localparam [5:0] p8 = (~&((!((&(2'd0))+(&(4'sd1))))||(((4'sd3)<(-2'sd0))/(3'sd0))));
  localparam signed [3:0] p9 = ((-4'sd7)!=(5'd2 * (~(~(2'd2)))));
  localparam signed [4:0] p10 = (5'd21);
  localparam signed [5:0] p11 = (-3'sd2);
  localparam [3:0] p12 = (2'd3);
  localparam [4:0] p13 = (((4'sd3)===(2'd2))/(2'd1));
  localparam [5:0] p14 = (~{({{(3'd3)}}>>>(~|((-3'sd2)?(5'd0):(3'sd2))))});
  localparam signed [3:0] p15 = ((~&((4'sd3)?(4'd7):(5'sd9)))?(|(-((2'sd0)%(-5'sd3)))):((~^(2'sd1))*((5'd4)%(2'd1))));
  localparam signed [4:0] p16 = {(-3'sd0)};
  localparam signed [5:0] p17 = (~(2'd3));

  assign y0 = {(-(-(p15?p14:p14))),((~p2)?(b3!==b4):(a1||p14)),(-((p5>=p3)+(a0===b5)))};
  assign y1 = (5'd29);
  assign y2 = (b1>>b1);
  assign y3 = (-5'sd1);
  assign y4 = {4{(^p9)}};
  assign y5 = (5'd3);
  assign y6 = {2{{2{$signed((a3^b0))}}}};
  assign y7 = (+({2{(!{4{p14}})}}?(|({2{p15}}&&(b4-b0))):(!((~a0)?(a2?p4:p6):(!p9)))));
  assign y8 = ((b5^~a4)?(a5?a1:a0):(~|a4));
  assign y9 = {4{$unsigned({1{(b3-b3)}})}};
  assign y10 = ((6'd2 * p1)-(b2||b5));
  assign y11 = (((b4>a1)^~{2{a4}})?((~^(&b1))>(&(&b0))):({3{b0}}|(a4?b1:b1)));
  assign y12 = ({{p4,p13},(p1>>>p4),{(~^p4)}}^(~&(~|{(a4===a3),(~&p13),(p1<<b2)})));
  assign y13 = (~^(~^((5'd7)>=(3'd7))));
  assign y14 = ((~|(+p14))<$signed((p12?p17:p6)));
  assign y15 = $signed({1{($signed(((p3|b5))))}});
  assign y16 = (~^{(&($unsigned((&$signed(((~^b5)))))))});
  assign y17 = ((p2?p13:p2)<={p7,p15,p13});
endmodule
