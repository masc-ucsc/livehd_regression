module expression_00575(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(!(&(|(4'd10))))}};
  localparam [4:0] p1 = (~&(-2'sd0));
  localparam [5:0] p2 = (-(5'd24));
  localparam signed [3:0] p3 = {{2{(3'd6)}},((3'sd2)?(-4'sd6):(3'd6))};
  localparam signed [4:0] p4 = (~{{((-2'sd1)<<(4'd8)),(!(5'd12)),(3'd6)},{((~(4'd7))>>>{(3'd5),(3'd5)})}});
  localparam signed [5:0] p5 = {{{{(-3'sd0),(5'sd0)}}},(((2'd3)!==(5'd19))?((5'd22)!=(5'sd10)):((2'd1)+(5'sd1)))};
  localparam [3:0] p6 = (~^((4'd10)<=(-3'sd3)));
  localparam [4:0] p7 = ((({2{(5'd15)}}!=((4'sd6)>(-2'sd1)))>>>({2{(2'd2)}}<{1{(3'd6)}}))!=={3{((5'sd4)&(-4'sd3))}});
  localparam [5:0] p8 = (|({((-2'sd0)===(2'd1)),((2'sd0)||(4'sd3)),((-3'sd2)-(2'd0))}>=(~&({(2'd0),(-4'sd6),(-5'sd5)}-(~|(2'sd1))))));
  localparam signed [3:0] p9 = (|(3'sd3));
  localparam signed [4:0] p10 = ((((-4'sd2)?(4'd11):(5'd5))&(((2'sd0)?(2'd2):(2'd3))^((2'd1)?(3'd3):(-2'sd0))))+(((-3'sd1)<(5'd11))?((2'd2)-(3'd1)):((4'd13)!==(2'sd1))));
  localparam signed [5:0] p11 = ((^{2{(-(4'd9))}})|({1{(-2'sd0)}}==={4{(4'sd6)}}));
  localparam [3:0] p12 = (((-2'sd1)/(4'd4))^~((2'd2)==(-4'sd3)));
  localparam [4:0] p13 = ((((-4'sd6)+(-2'sd1))||(-5'sd11))>=(3'sd3));
  localparam [5:0] p14 = {((2'd2)?(-2'sd1):(5'd10)),{3{(-3'sd3)}}};
  localparam signed [3:0] p15 = (((3'd4)>(2'sd1))===((4'sd0)+(5'sd15)));
  localparam signed [4:0] p16 = (2'sd0);
  localparam signed [5:0] p17 = (((((5'd7)<<(4'd1))>=((4'd11)!==(2'd3)))<{1{{2{(5'd11)}}}})&&(|(((4'sd7)<(-3'sd2))==={2{(2'd1)}})));

  assign y0 = (-4'sd7);
  assign y1 = (((~^{1{(|(|{4{p9}}))}}))<=(+(|(!$signed((b2^b0))))));
  assign y2 = ((p11>=p7)<<<(a5+a0));
  assign y3 = (-2'sd0);
  assign y4 = ($unsigned(((b3!==a0)))<<<$unsigned(((b2!==a0)>=(4'sd1))));
  assign y5 = (a5?p16:a0);
  assign y6 = (-(3'sd0));
  assign y7 = (((p12?p3:a2)||(+b5))^{(+b2),(p5?p5:p13)});
  assign y8 = (5'd21);
  assign y9 = ((((~&b2)||(b3&&a1))+(3'd3))!==(-3'sd1));
  assign y10 = (a4<<p0);
  assign y11 = ((2'd0)==((^$unsigned(p17))?(-5'sd9):(b3?p12:p0)));
  assign y12 = {2{{1{{{1{b2}},{3{p1}},{2{b2}}}}}}};
  assign y13 = ($unsigned((-(-((~(b3?p11:a3))!={(-$unsigned((~a4)))})))));
  assign y14 = ((~(~(4'd2 * (b1?b0:a2))))||(~|(!((&(a0?b1:a5))&&(&(b0>=a4))))));
  assign y15 = ((^({1{p14}}>>{3{p17}}))^(2'd3));
  assign y16 = (3'sd1);
  assign y17 = (3'd7);
endmodule
