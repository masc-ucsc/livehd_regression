module expression_00116(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(+((4'd12)+(5'd19)))}};
  localparam [4:0] p1 = ((3'sd0)^~(-4'sd4));
  localparam [5:0] p2 = (-2'sd0);
  localparam signed [3:0] p3 = (((-2'sd1)<(3'd1))<=((5'd22)?(4'd6):(2'd0)));
  localparam signed [4:0] p4 = {{(5'd2 * (2'd3)),((5'd24)+(2'd2)),{(2'd1),(5'd21),(-2'sd1)}},(6'd2 * {((2'd2)<=(2'd2))})};
  localparam signed [5:0] p5 = ((4'd1)?(4'sd0):(-3'sd3));
  localparam [3:0] p6 = (((4'd8)?(5'sd4):(5'sd7))<((5'd19)!=(2'sd1)));
  localparam [4:0] p7 = (4'd13);
  localparam [5:0] p8 = ((((-4'sd1)==(-3'sd2))<=(-(3'd0)))?((4'd10)<=((5'sd14)?(5'd24):(4'd3))):(2'd3));
  localparam signed [3:0] p9 = ((((5'd31)?(-2'sd1):(4'd12))<{1{(2'd2)}})?(((5'd12)===(4'd3))+((3'd0)^(3'sd0))):(((-3'sd0)||(5'd0))?{4{(2'sd1)}}:((3'sd0)?(3'd4):(4'sd2))));
  localparam signed [4:0] p10 = (~|(3'd7));
  localparam signed [5:0] p11 = (|((|({3{(3'sd2)}}&&((4'sd6)^(5'd10))))>{4{(4'sd4)}}));
  localparam [3:0] p12 = ((~|((-5'sd7)?(5'd0):(-3'sd2)))?(((4'sd4)!==(-4'sd2))^((3'd6)<(5'd7))):(+((5'sd3)?(2'd2):(5'sd11))));
  localparam [4:0] p13 = (-2'sd0);
  localparam [5:0] p14 = (|(-2'sd0));
  localparam signed [3:0] p15 = {2{(2'sd1)}};
  localparam signed [4:0] p16 = {(~^(^(^(~&{(4'd4)})))),{(|(3'sd3)),(&(4'd4)),{(3'd6)}}};
  localparam signed [5:0] p17 = ((~^(4'sd1))<<<((2'sd0)?(5'sd8):(4'sd3)));

  assign y0 = (-2'sd0);
  assign y1 = ((6'd2 * $unsigned((p5>>p17)))>(4'sd5));
  assign y2 = {$signed({$unsigned({(~p3),(+p11)}),($signed($signed({b2,b2,p7})))})};
  assign y3 = ((^((!(p9?p0:p9))|(p9?a1:p5)))!=(((|b0)?(p7&&p9):(b1?p15:p11))>>>((!p8)?(p12^p9):(p12?p15:p1))));
  assign y4 = (&(((a2/b5)||(b5&&p9))|((b3?p14:p8)?(a5?b5:b2):(p11/a5))));
  assign y5 = (-4'sd2);
  assign y6 = (~(~|a0));
  assign y7 = ({4{a3}}?(a4):(+a4));
  assign y8 = $unsigned({{p1}});
  assign y9 = ({1{{3{(|{1{p9}})}}}});
  assign y10 = ((b2?a5:p9)/b2);
  assign y11 = (~&$unsigned(b0));
  assign y12 = $signed((4'd2 * (a2>b1)));
  assign y13 = {4{((p10<<<p5)<<<(p0&&p6))}};
  assign y14 = {1{(($signed(a1)?(b2?b0:b2):(a3^~a5))!==(!{1{({4{a0}}<<(b0?a2:a5))}}))}};
  assign y15 = (6'd2 * (b0!=p6));
  assign y16 = {{1{(!(~{4{b1}}))}},{$signed({{1{b3}}}),{4{b3}}}};
  assign y17 = ({(5'd2 * p13),{3{a5}},(a5===b5)}&&(((p10&p4)-(p12?a0:a2))>{{p2},{1{p0}},(p2?b1:p9)}));
endmodule
