module expression_00929(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(|{3{((5'd18)?(-3'sd1):(2'sd0))}}));
  localparam [4:0] p1 = {4{((-3'sd2)?(2'd0):(2'd0))}};
  localparam [5:0] p2 = ((|(((5'd6)|(2'd1))^(~|(5'd28))))>(((-2'sd0)===(2'd0))&&(^(4'd6))));
  localparam signed [3:0] p3 = {(4'd13),(2'd0)};
  localparam signed [4:0] p4 = (((5'd8)/(5'd0))?(6'd2 * (3'd6)):(~((-2'sd0)?(5'd26):(4'sd5))));
  localparam signed [5:0] p5 = (4'd0);
  localparam [3:0] p6 = (3'd0);
  localparam [4:0] p7 = (({(4'sd1),(-2'sd1),(2'd1)}?(|(2'sd0)):{(-5'sd14),(3'sd3),(2'sd1)})<<<(^(((5'd12)==(-5'sd8))!=(~|(3'd2)))));
  localparam [5:0] p8 = (5'd2 * (2'd0));
  localparam signed [3:0] p9 = {3{((4'd7)!==(4'sd3))}};
  localparam signed [4:0] p10 = (2'd0);
  localparam signed [5:0] p11 = ((~((4'd11)>>(3'd3)))+(3'd5));
  localparam [3:0] p12 = (+((((4'sd1)<<(2'sd1))>((5'd13)-(-4'sd4)))<<<{((2'd3)!=(2'd3)),(6'd2 * (5'd18)),((3'sd3)&(-2'sd1))}));
  localparam [4:0] p13 = (&{(~^(2'sd1)),(~&(^{(3'd4),(2'd3),(4'd9)})),(-(3'd2))});
  localparam [5:0] p14 = (-2'sd0);
  localparam signed [3:0] p15 = (~(3'd7));
  localparam signed [4:0] p16 = ((2'sd0)>{(5'd5),(5'sd13),(2'd3)});
  localparam signed [5:0] p17 = (-(-2'sd1));

  assign y0 = (((p7?p0:p2)<<<(~(-p13)))?(~|(^{2{{4{a0}}}})):((p15?a4:a1)?(-5'sd8):(&b0)));
  assign y1 = (~&($signed(p7)?(!p6):(p1||p16)));
  assign y2 = (((p4-p10)^(p2&a4))?{(p9<p5),{p15,b5,a2}}:(4'sd5));
  assign y3 = (+(((-p4)+(p11||p8))>>>((!p10)<<(p1-p0))));
  assign y4 = (~^(|(p2>>a4)));
  assign y5 = {(!((p3>>b3)+{p14,b0,p16})),(!((p7!=p2)>={a5,p15}))};
  assign y6 = (p15&&p7);
  assign y7 = (3'd3);
  assign y8 = (((p15?p3:p17)==(p16?p10:p0))?((p2!=p16)=={(4'd2 * p1)}):({p3,b3,p8}^~{p13,p1,p6}));
  assign y9 = {4{(~|{p11,p2})}};
  assign y10 = {b0,p3,b5};
  assign y11 = {4{(^p7)}};
  assign y12 = (((b0===a3)<{4{p15}})||(4'd2 * (a0>>b1)));
  assign y13 = ((+{4{b5}})?(~^(b2^~a0)):{3{a0}});
  assign y14 = {4{{4{a3}}}};
  assign y15 = (~(~^(5'd2 * (4'd12))));
  assign y16 = $unsigned($signed(($unsigned((p9?p3:p4))&&(p1?p6:b5))));
  assign y17 = (-((~^{{1{p3}},(p6?b1:b2)})^~(2'd0)));
endmodule
