module expression_00982(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{{(3'd3)}},{(-4'sd3),(2'd2),(5'd23)},{{(4'd10),(4'd10),(-5'sd13)}}};
  localparam [4:0] p1 = (+(~&(&{(~|{(4'd3),(2'sd0),(4'd9)}),{(~^(5'd22))}})));
  localparam [5:0] p2 = ((((-3'sd0)<(2'sd1))>>((-4'sd7)*(4'd14)))<<(((-3'sd3)>(5'd4))==((-5'sd6)<=(4'd14))));
  localparam signed [3:0] p3 = (5'd23);
  localparam signed [4:0] p4 = (!((^(4'd2))===((-3'sd3)?(-4'sd4):(2'd0))));
  localparam signed [5:0] p5 = ({(3'sd1)}?((2'd0)>=(-4'sd6)):((5'd0)===(-4'sd0)));
  localparam [3:0] p6 = ({2{((4'd0)<<<(4'd9))}}||(2'sd1));
  localparam [4:0] p7 = (|{(-4'sd1),(-(-2'sd0))});
  localparam [5:0] p8 = ((((2'd3)+(3'd7))?((-2'sd1)?(4'd4):(2'sd1)):((5'd19)<<<(2'd2)))==(((-5'sd2)?(3'd7):(5'd27))?((3'd2)+(4'sd3)):{(5'sd9),(3'd7),(3'd0)}));
  localparam signed [3:0] p9 = (~(|(~&((+((-4'sd6)>(2'sd0)))>(~((2'sd0)<=(3'd6)))))));
  localparam signed [4:0] p10 = ((&((5'sd14)<=(5'd1)))-((5'd21)===(3'd5)));
  localparam signed [5:0] p11 = ({((-4'sd6)&(2'd3)),(&(4'd2))}?(+(4'd10)):(((-3'sd1)?(2'd0):(-4'sd0))?(4'sd2):(~&(4'sd1))));
  localparam [3:0] p12 = {{1{{(-3'sd0),(-4'sd6),(5'sd2)}}},((-2'sd1)?(3'd7):((-3'sd2)>>>(5'd24))),(5'sd14)};
  localparam [4:0] p13 = ({{(-5'sd2),(3'd7)},{2{(4'd2)}},(~|(4'd2 * (4'd4)))}<=(((3'd7)?(2'sd0):(2'd2))^~((2'd2)?(5'd12):(4'sd0))));
  localparam [5:0] p14 = ((2'd0)||(2'sd1));
  localparam signed [3:0] p15 = ((((-3'sd2)?(3'sd1):(-3'sd0))?((-4'sd0)<<(4'd1)):((4'd2)?(4'd15):(2'sd1)))&&(((3'sd1)?(3'd0):(5'd2))^((5'd5)||(2'd0))));
  localparam signed [4:0] p16 = ((^(3'd5))?((3'd7)?(4'd4):(5'd10)):(-(3'sd3)));
  localparam signed [5:0] p17 = (((3'd2)?(4'd3):(3'sd1))?((5'sd6)?(-5'sd15):(3'd7)):(^{(5'd22)}));

  assign y0 = ((p10?b5:p15)>(b4?a1:a4));
  assign y1 = ((b0?a1:b0)!==(b2?b0:a4));
  assign y2 = (|(p10>>p0));
  assign y3 = {4{((a1!==b3)<=(a0^a2))}};
  assign y4 = (4'd11);
  assign y5 = ((p12&b5)<<<{a2,b2});
  assign y6 = (-(b3===b5));
  assign y7 = ((5'sd14)&(^(p4&&a5)));
  assign y8 = ({(a3?a0:a5),{p16,b0},{b3}}?((a4>>a2)!==(a4?a3:a4)):{(b5+a3),(p17>b4)});
  assign y9 = ({(~&{a0,p7})}<=(+((~|{b2,b1}))));
  assign y10 = (({1{(p15^p17)}}>>>{{p11,p5,p6}})^~{{2{{3{p7}}}},{4{p5}}});
  assign y11 = {3{{2{{2{a1}}}}}};
  assign y12 = (|(-(((p10>>p0)<<<(~&a1))+(~&(|(&p2))))));
  assign y13 = ({{(a4!==a0)}}<((b2!==a0)&&{a2,a1,b1}));
  assign y14 = {3{(a5+a2)}};
  assign y15 = {b3,p15,b1};
  assign y16 = {2{((!(p8!=p7))&&((!p1)+{3{p0}}))}};
  assign y17 = (|$unsigned(((p7?p12:p10)?$unsigned(b0):(p13))));
endmodule
