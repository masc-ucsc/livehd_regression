module expression_00596(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^((2'sd0)!==(4'd9)))*((-3'sd1)?(5'd28):(-4'sd0)));
  localparam [4:0] p1 = (((3'd5)!==(4'd15))?((2'd0)-(-3'sd3)):((5'd28)?(3'd1):(4'sd6)));
  localparam [5:0] p2 = (((4'd0)^~(3'd1))/(2'd2));
  localparam signed [3:0] p3 = (5'sd15);
  localparam signed [4:0] p4 = ((-(~^{2{{3{(5'd31)}}}}))+(~&(((5'd0)!=(-2'sd1))||((3'd6)!=(-2'sd0)))));
  localparam signed [5:0] p5 = (~&(+{1{(~(&({1{((!(4'd12))<<<{2{(2'd3)}})}}&&{4{(-2'sd0)}})))}}));
  localparam [3:0] p6 = {(((2'd0)?(2'sd0):(2'sd0))!==((-2'sd1)^~(-2'sd0)))};
  localparam [4:0] p7 = (-2'sd0);
  localparam [5:0] p8 = ((-3'sd2)===(5'd23));
  localparam signed [3:0] p9 = ((3'd3)+(4'd12));
  localparam signed [4:0] p10 = (~&{3{(~&(((4'd13)&&(5'd16))<<((2'd3)||(5'd23))))}});
  localparam signed [5:0] p11 = (((-2'sd0)&(5'd2))/(4'd4));
  localparam [3:0] p12 = ({1{{1{(((4'd12)!=(3'sd0))<(!(2'd2)))}}}}>>(+(((5'd30)|(5'd18))>((-2'sd0)?(5'd10):(2'd0)))));
  localparam [4:0] p13 = ((4'd15)?(-3'sd2):(-3'sd2));
  localparam [5:0] p14 = ({{(^(5'd26)),{(5'd11)}}}&(((2'd3)===(3'sd1))===(+(3'd5))));
  localparam signed [3:0] p15 = (((3'd0)<(2'sd1))&&((4'sd7)!=(5'd5)));
  localparam signed [4:0] p16 = (~|(^{(((4'd3)&(2'd3))?{3{(5'sd14)}}:((3'd4)?(2'd3):(3'd7))),(5'sd11)}));
  localparam signed [5:0] p17 = (((~&(5'd14))>=((3'd3)&(3'd4)))<<<(~((5'sd10)?(4'sd4):(4'd13))));

  assign y0 = (^(4'sd0));
  assign y1 = (((~|(+b1))*(~(b5<=a0)))<<(^(2'd1)));
  assign y2 = ((b1<=p10)^$unsigned(b0));
  assign y3 = ((-5'sd14)-(2'd3));
  assign y4 = (((-3'sd2)>(p17<<b1))>>$signed((4'd3)));
  assign y5 = (2'sd1);
  assign y6 = (((a4<<<a0)?(~&(~|a0)):(!(b0===a5)))!==((6'd2 * a1)?$signed((a3?a2:a1)):$unsigned((b2===b3))));
  assign y7 = {4{{2{(a2!=a4)}}}};
  assign y8 = (|{2{{(p4?p5:p10)}}});
  assign y9 = (4'd2);
  assign y10 = ({2{(+(~(p9&a3)))}}+(((p1<<p2)==(!p0))>={1{(p15!=p8)}}));
  assign y11 = ({1{b0}}?{3{p9}}:{1{b0}});
  assign y12 = ({4{a5}}||(^(~|(-p11))));
  assign y13 = (~|{(3'd0),(p11?b5:b1),(4'd14)});
  assign y14 = (4'd0);
  assign y15 = {(~(3'sd3)),(~^{(4'd9)}),({(a2>=a4)}-(b4!==a0))};
  assign y16 = (+a5);
  assign y17 = (3'sd3);
endmodule
