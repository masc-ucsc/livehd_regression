module expression_00014(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^{(+(&{(2'sd0),(3'sd2)}))})!==(&(((2'd3)<<<(2'sd1))+{(-(4'd8))})));
  localparam [4:0] p1 = (+(-3'sd2));
  localparam [5:0] p2 = (~|(~|(~&(|(~|(&(|(+(5'd16)))))))));
  localparam signed [3:0] p3 = {3{{(-5'sd1),(-2'sd0)}}};
  localparam signed [4:0] p4 = (~|(5'd28));
  localparam signed [5:0] p5 = (-2'sd1);
  localparam [3:0] p6 = {{(+(5'd21))},{4{(-5'sd6)}},(6'd2 * (4'd5))};
  localparam [4:0] p7 = (5'd25);
  localparam [5:0] p8 = (+(-2'sd1));
  localparam signed [3:0] p9 = (({1{((2'd0)-(-5'sd4))}}^{3{(3'sd2)}})<<(((5'sd11)<<<(-2'sd1))<<<((4'sd6)>>>(-3'sd2))));
  localparam signed [4:0] p10 = (~&(~((3'sd0)<=(4'sd2))));
  localparam signed [5:0] p11 = ({4{(2'd1)}}-(~^((2'd3)<(3'sd3))));
  localparam [3:0] p12 = (3'd0);
  localparam [4:0] p13 = (~&(-3'sd1));
  localparam [5:0] p14 = {1{(5'd8)}};
  localparam signed [3:0] p15 = ((~^(&((3'd4)|(-5'sd3))))?((-4'sd5)?(-5'sd6):(-3'sd3)):{3{(2'd1)}});
  localparam signed [4:0] p16 = {4{(2'd1)}};
  localparam signed [5:0] p17 = ({1{({1{(3'sd1)}}!={(-5'sd2),(5'd30)})}}<={((4'sd6)^~(2'd1)),((4'sd4)<<(-3'sd3)),((5'd24)+(4'd15))});

  assign y0 = {3{(&p9)}};
  assign y1 = $unsigned({(&((~((b3)))<=(a1?b3:b5))),{(-(b2+a3)),(|(^{b2,a2,a0}))}});
  assign y2 = {(-5'sd2),(~{a1})};
  assign y3 = (^({p11,a1,p15}?(p1>>p7):$unsigned(p13)));
  assign y4 = (5'd4);
  assign y5 = (~&((-(!(-a2)))?(^(~|(p5>>>a2))):((~^p12)*(-3'sd3))));
  assign y6 = (($signed((~^((-4'sd6)<<<(!p14)))))-(|{(5'd16),(|a3),(~p3)}));
  assign y7 = (((a1?b5:b2)!=={b3,b2,b4})==((!b3)?(-5'sd14):(a4|a3)));
  assign y8 = {3{(p12?p16:p3)}};
  assign y9 = ({3{(p11<<<a5)}}-{1{((p11^~b0)^{2{p9}})}});
  assign y10 = (({4{a5}}=={{{b0,p4}}})<={2{{(p3?a5:p11),{4{a2}}}}});
  assign y11 = ((-5'sd1)>$unsigned((~((~(a2|p0))>>>$unsigned((b4||b5))))));
  assign y12 = (5'd10);
  assign y13 = {{{(b4<<p10)},(({4{b3}}))}};
  assign y14 = (p9<=p6);
  assign y15 = (2'd2);
  assign y16 = {((a2!==a1)?(p15>p9):(b2<<p2)),((p10<a4)>>{a1,b4})};
  assign y17 = (((5'd26)<<(-3'sd0))&&(4'd10));
endmodule
