module expression_00486(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(3'd5));
  localparam [4:0] p1 = ((&((~^(2'sd1))?(|(3'd2)):((-5'sd6)^~(4'd4))))&&(((4'sd3)^~(3'd2))?((5'sd12)<=(-3'sd1)):((5'sd10)?(2'sd1):(4'sd4))));
  localparam [5:0] p2 = (^(-2'sd1));
  localparam signed [3:0] p3 = {(~|({(2'd0),(5'd22),(3'sd1)}?{3{(5'd20)}}:((3'd1)?(2'd1):(5'd13)))),(-4'sd0)};
  localparam signed [4:0] p4 = {1{{2{(~&((3'd4)?(4'd13):(4'd1)))}}}};
  localparam signed [5:0] p5 = (~&((~|((-(2'sd0))*(-(4'd4))))?(~&(((-4'sd6)+(2'sd1))&((-3'sd1)-(5'd11)))):((4'd2 * (3'd3))&&((-3'sd3)||(4'd13)))));
  localparam [3:0] p6 = (~|((~|(5'sd12))?(^(|(4'd10))):((4'd8)?(-4'sd5):(2'd0))));
  localparam [4:0] p7 = ((-5'sd12)-(-2'sd1));
  localparam [5:0] p8 = (~(2'd2));
  localparam signed [3:0] p9 = (!((~|((-5'sd1)?(5'd20):(-2'sd0)))?((2'd1)?(3'sd0):(-4'sd0)):(+(&(4'd15)))));
  localparam signed [4:0] p10 = (~^((^((|(3'd3))>>>((-2'sd0)==(-3'sd1))))!==((-(~&(5'sd11)))==(~^(~^(4'd8))))));
  localparam signed [5:0] p11 = (+(5'sd11));
  localparam [3:0] p12 = (3'd3);
  localparam [4:0] p13 = (((4'd13)?(5'd18):(5'd11))?((5'd7)?(-2'sd0):(2'd0)):((3'sd0)?(3'sd0):(4'd7)));
  localparam [5:0] p14 = (-2'sd0);
  localparam signed [3:0] p15 = ((|(-3'sd0))===(-(-3'sd1)));
  localparam signed [4:0] p16 = (~(2'd2));
  localparam signed [5:0] p17 = {4{(2'sd1)}};

  assign y0 = (2'd1);
  assign y1 = {{p9},(-p15),(a3?b5:b3)};
  assign y2 = ((&(-$unsigned(((2'd1)>>>(p6>=p16)))))>>(-2'sd1));
  assign y3 = (~^(({2{p5}}?{4{p0}}:{3{b3}})!={2{((p5>b5)-(p12&&p17))}}));
  assign y4 = (3'sd0);
  assign y5 = (a0<=a3);
  assign y6 = (^({2{p9}}|(a2!==a4)));
  assign y7 = {2{((a3?p4:a0)-(p10<<<a4))}};
  assign y8 = (~(+(-4'sd0)));
  assign y9 = (^((~(p12||b2))?((p1>b2)!=(b2===b1)):((~a0)<=(~|b2))));
  assign y10 = (&({2{a3}}===(a1?b2:b5)));
  assign y11 = (!{3{{1{b5}}}});
  assign y12 = {({(-4'sd2),$signed(b4)}>(3'sd1)),(3'sd1)};
  assign y13 = ({2{({1{p7}})}}?(3'd1):(-(^(|{2{p12}}))));
  assign y14 = ((b3?b2:b2)!=((b4==b0)/a4));
  assign y15 = {4{p7}};
  assign y16 = (5'sd12);
  assign y17 = ((2'd1)+(a3>>>a5));
endmodule
