module expression_00961(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(~&(2'sd0)),((-2'sd0)?(-3'sd1):(5'sd5))}?({(3'sd1)}?{(4'd5)}:(+(5'd19))):((+(4'd12))?(~(-2'sd1)):((5'd23)?(5'sd1):(-4'sd0))));
  localparam [4:0] p1 = {(|(-4'sd6))};
  localparam [5:0] p2 = (-5'sd3);
  localparam signed [3:0] p3 = (&((~|(4'd2 * (!(!(4'd12)))))!==((5'd2 * (2'd3))!=((4'd11)-(-5'sd8)))));
  localparam signed [4:0] p4 = ((((-2'sd0)?(5'd30):(-5'sd5))?((4'd11)?(2'd1):(-3'sd1)):((2'd3)&&(-4'sd5)))^~(6'd2 * {2{(5'd2)}}));
  localparam signed [5:0] p5 = (&{2{{{1{((4'd5)===(-4'sd5))}}}}});
  localparam [3:0] p6 = (5'd7);
  localparam [4:0] p7 = (~&{(2'sd0),(4'd0),(5'd21)});
  localparam [5:0] p8 = (!((-((5'd4)^(-5'sd1)))>((^(4'd12))|(&(2'sd0)))));
  localparam signed [3:0] p9 = (&(&(4'sd3)));
  localparam signed [4:0] p10 = (~|{4{(4'sd5)}});
  localparam signed [5:0] p11 = (+({4{((-4'sd5)!==(5'sd7))}}>>((~(~|(-4'sd4)))===((4'sd0)?(4'd8):(-5'sd10)))));
  localparam [3:0] p12 = (((2'd1)?(4'd12):(5'd5))&&((2'd1)?(4'd7):(-2'sd0)));
  localparam [4:0] p13 = (&((+((3'd1)-(5'd15)))+((4'd1)^(5'd14))));
  localparam [5:0] p14 = {{(((2'sd1)&(4'sd1))==((5'sd3)>(5'sd9))),(((4'sd7)?(-2'sd1):(5'd22))=={(4'd15)}),{((4'd13)&(-3'sd0)),(6'd2 * (5'd31)),((-4'sd3)!=(-3'sd3))}}};
  localparam signed [3:0] p15 = {(!(2'sd0)),((-5'sd11)?(5'd3):(5'd18))};
  localparam signed [4:0] p16 = (&(^(((3'd0)>>(3'd3))-((2'd1)|(-2'sd1)))));
  localparam signed [5:0] p17 = {{(5'sd13),(-4'sd2),(2'd0)},({(4'd12)}|(-(3'd0))),{(2'd1),(4'sd1),(2'd0)}};

  assign y0 = (b4?a4:b2);
  assign y1 = ((b1?a5:p2)?(a2?p17:a3):(p15&&b2));
  assign y2 = {{(~^p9),{a1,a0,p16}},(&((a2||p13)>=(3'sd3)))};
  assign y3 = (({p0,b2,a3}?(!b5):(2'd1))?((5'd29)?(-b4):(~b2)):(&{(a5?b5:b3),(^b2)}));
  assign y4 = (~(3'sd0));
  assign y5 = (((~|p8)?(p1?p1:p14):(b4===b1))||(~|(p2?p16:p3)));
  assign y6 = ((({a0}||(a3!==a4))<=({3{p16}}>>>(p12^~a2)))^~{{{4{b5}}},(b3<b0),{4{b4}}});
  assign y7 = ({a3,a3,a5}===(4'd1));
  assign y8 = (|(+p5));
  assign y9 = ((-((b1&b2)<<{(a4?b0:a1)}))|((b2<p4)?{(p15>>a2)}:(b3^~b0)));
  assign y10 = $signed({{{{b3,a2,a0}}},$unsigned($unsigned($unsigned({b2,b4}))),{{{a3,a4}}}});
  assign y11 = ((&(^(($signed(((-$signed((b4<<b4)))))&&((|(a1>b5))-$unsigned((|a4))))))));
  assign y12 = (((b1?a1:a0)/p16)?((a0===b0)?(+a4):(p9&p17)):(~(~^(-(p9?b3:p11)))));
  assign y13 = (^{{(p11&&p15)}});
  assign y14 = ((a2>=p5)?(+(3'd1)):(~|(p5?p8:p2)));
  assign y15 = (!((-2'sd0)?{p16}:(~&p9)));
  assign y16 = ((|(5'sd13))>(-({(a2^a5)}?(5'd17):(-(-4'sd6)))));
  assign y17 = ((p14==p0)?(-(&a3)):(p14^~p0));
endmodule
