module expression_00224(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd12)|{(~^(~(5'd1))),((5'd25)>(-2'sd0))});
  localparam [4:0] p1 = {(~&((3'sd1)<=(3'd6))),{(-4'sd5),(3'd7),(-3'sd0)},((3'd7)&(5'd2))};
  localparam [5:0] p2 = ((3'd5)!=(2'sd1));
  localparam signed [3:0] p3 = {(((-5'sd0)-(5'd3))>>>((3'd4)!==(3'd6))),(4'd2 * (4'd9)),(~(((2'sd0)==(3'd4))||(-4'sd7)))};
  localparam signed [4:0] p4 = ((4'd2 * {2{(5'd26)}})|{2{((2'd3)|(3'd2))}});
  localparam signed [5:0] p5 = (-({1{(-{1{(4'd6)}})}}?((-2'sd0)?(5'sd2):(5'd11)):(^(3'sd2))));
  localparam [3:0] p6 = (-(-4'sd4));
  localparam [4:0] p7 = (~^{4{{3{(-3'sd0)}}}});
  localparam [5:0] p8 = (|(|(&({((3'd7)^~(4'd12)),((4'd4)!=(-3'sd0)),{(3'sd2),(4'd3),(3'd6)}}||((5'sd15)^~{(2'd2),(-2'sd0)})))));
  localparam signed [3:0] p9 = (~|(-2'sd0));
  localparam signed [4:0] p10 = ((-3'sd2)<<<(4'd1));
  localparam signed [5:0] p11 = (((4'sd3)^(4'd0))?((2'd2)>>(5'sd3)):((-3'sd1)?(4'd0):(2'sd0)));
  localparam [3:0] p12 = (~^(|(&((2'sd0)?(2'd2):(5'sd5)))));
  localparam [4:0] p13 = (|(~&(|{((2'sd1)?(-4'sd7):(2'd2))})));
  localparam [5:0] p14 = {4{{(-3'sd2),(-4'sd3),(-5'sd7)}}};
  localparam signed [3:0] p15 = {1{(^((4'd8)||(5'd22)))}};
  localparam signed [4:0] p16 = ({2{{(2'd0)}}}&&{((4'd13)?(-2'sd1):(2'd2)),((2'sd0)!==(4'sd1))});
  localparam signed [5:0] p17 = ((-4'sd3)?(4'd3):(2'd3));

  assign y0 = (b3?b4:p17);
  assign y1 = (^{b5,p17,b4});
  assign y2 = $unsigned((^((+((a0<=p6)!=(p5?p14:b4)))>>(~(+((p6?p4:a2)?(p2<<<p5):(p9>=p11)))))));
  assign y3 = ((p3)?(+b3):(^b4));
  assign y4 = (&(-2'sd0));
  assign y5 = (&(((-(+p10))+(|(~|p15)))||((-(~^b4))!==(~(+b1)))));
  assign y6 = ((b0*p14)?(a0?p2:a3):$signed(a3));
  assign y7 = ({2{{2{p8}}}}?{2{(p9?a5:p9)}}:({1{p17}}?(p15?p5:a0):(p4?p15:p15)));
  assign y8 = (~{(&((p12+p15)-{(|p3)}))});
  assign y9 = (+(!(3'd7)));
  assign y10 = ((!{1{(~^({2{a5}}?{1{p4}}:(a5?b3:b0)))}})|(({b5,a0,b3}&(~^a4))<<((a0?p4:a4)&&(|p4))));
  assign y11 = ((~|($unsigned((p2>>p1))+(!(~^(b4>>a1)))))&(+$unsigned({{p12,b1,b3},(b5&p6),(!(a2>>b3))})));
  assign y12 = ((~^(p5?p8:p2))?(p11?p4:p6):(p5?p7:p16));
  assign y13 = ({2{(a2-p14)}}-({1{(p8>>b0)}}<{3{p2}}));
  assign y14 = {$signed((+(~^p8))),((p0!=p3)==(3'd5))};
  assign y15 = {2{{(a4>>>p7)}}};
  assign y16 = (4'd10);
  assign y17 = (+$unsigned(a2));
endmodule
