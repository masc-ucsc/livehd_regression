module expression_00154(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({4{(3'd7)}}<<{(-5'sd12)})?{((5'd8)>>(2'd1)),{(5'd9)}}:((3'd2)?(4'd15):(-5'sd14)));
  localparam [4:0] p1 = (6'd2 * ((5'd1)&&(2'd3)));
  localparam [5:0] p2 = (+(2'd0));
  localparam signed [3:0] p3 = {3{((4'd2 * (4'd9))|(4'd6))}};
  localparam signed [4:0] p4 = (+(-2'sd0));
  localparam signed [5:0] p5 = (4'sd4);
  localparam [3:0] p6 = (&((-4'sd3)===(^((4'sd7)<<<(4'd4)))));
  localparam [4:0] p7 = (3'd4);
  localparam [5:0] p8 = (6'd2 * ((3'd1)>>>(4'd10)));
  localparam signed [3:0] p9 = (((4'd7)<=(2'sd1))?(5'sd6):(5'sd15));
  localparam signed [4:0] p10 = ((~&(~|(!({4{(2'sd0)}}>={(3'd5),(2'd3),(-4'sd2)}))))-((~{1{(-3'sd1)}})<<<(2'd3)));
  localparam signed [5:0] p11 = {4{(-3'sd3)}};
  localparam [3:0] p12 = (^({(~(~&{(4'sd0)}))}?{(~^(2'd3)),((-5'sd7)?(4'd5):(-3'sd2))}:(-(!(&((5'd16)>>>(2'sd1)))))));
  localparam [4:0] p13 = (+(4'd2 * (4'd6)));
  localparam [5:0] p14 = (~{4{((5'd30)>>(4'sd2))}});
  localparam signed [3:0] p15 = ((2'd0)<<<(5'd13));
  localparam signed [4:0] p16 = (~&((3'd5)==(5'd6)));
  localparam signed [5:0] p17 = (((2'd2)|(3'sd3))!=(3'd2));

  assign y0 = ({3{(3'd7)}}^{4{{1{p2}}}});
  assign y1 = (((2'd2))|{((5'sd3)-(2'd2))});
  assign y2 = ({{1{a2}},(a3!==b1),(p4?a0:p16)}^~((p16?a0:b0)!=(p15?b5:a2)));
  assign y3 = (((-2'sd1)>=((3'sd3)||(-b4)))>=(5'd23));
  assign y4 = ((&{{b5,a2,a2},(b5<=a4)})==={3{(a0||b0)}});
  assign y5 = (a1|b2);
  assign y6 = ((5'd31)&&({p12,p9,p11}>=(b1||p12)));
  assign y7 = (|(~&p11));
  assign y8 = (({a4,b4,p12}&((b1<<<b0))));
  assign y9 = {4{b1}};
  assign y10 = (&{{1{{2{{4{(p15^~p14)}}}}}}});
  assign y11 = (((a3^a4)==(a4==b5))===(&(b5+a4)));
  assign y12 = {b2,p12};
  assign y13 = ((p6?a1:p15)<=(p5?p11:p16));
  assign y14 = (~{(~{(-a5),(~|b4),(!a4)}),(|{{b2,b2},(+{a4,a3,a5})})});
  assign y15 = (p7?a0:p11);
  assign y16 = ($signed((5'd6))<=(~^(2'd2)));
  assign y17 = ((4'd12)?$unsigned((4'd11)):((-3'sd2)?(2'sd1):(b0!==b0)));
endmodule
