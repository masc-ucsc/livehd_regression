module expression_00304(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({(5'd14)}>(~(5'sd0)))>>>(-((5'sd10)?(4'd7):(3'd5))));
  localparam [4:0] p1 = (+((~|(-(-4'sd4)))+(~(-5'sd10))));
  localparam [5:0] p2 = ((-2'sd0)?(3'sd0):(2'd1));
  localparam signed [3:0] p3 = ((^(((4'd0)?(3'sd0):(3'd2))^{3{(-4'sd5)}}))=={4{{3{(5'd24)}}}});
  localparam signed [4:0] p4 = ((5'd15)^(4'd9));
  localparam signed [5:0] p5 = ((((-5'sd11)<<<(-3'sd1))&&((2'sd1)!==(5'sd2)))&(((5'sd9)^~(5'd0))<<(!(4'd2 * (2'd3)))));
  localparam [3:0] p6 = (-{(~^{(~(4'd15)),{2{(-3'sd3)}}}),{(&(2'sd1)),{(2'd2),(2'd1),(2'd0)},{(4'd14),(3'sd3)}},(&{{(-2'sd1),(-5'sd10)},{(-5'sd13),(4'd12),(5'd19)}})});
  localparam [4:0] p7 = {2{(~^(~^((4'd2)?(2'd2):(5'sd4))))}};
  localparam [5:0] p8 = ((5'd20)<<<((2'sd1)+((2'sd0)<=(2'sd0))));
  localparam signed [3:0] p9 = ((-5'sd10)>{(-4'sd4),(2'sd0),(-2'sd1)});
  localparam signed [4:0] p10 = (|({(4'sd1),(2'd2),(-2'sd0)}^~((5'sd7)>=(5'sd15))));
  localparam signed [5:0] p11 = {(3'd0),(5'd10),(5'd7)};
  localparam [3:0] p12 = (&{(5'd15),{(~|(5'd19)),(5'd30),{(2'd2)}}});
  localparam [4:0] p13 = (3'sd0);
  localparam [5:0] p14 = (6'd2 * (|((4'd15)<(3'd1))));
  localparam signed [3:0] p15 = {2{({1{(2'd1)}}?((2'd1)<(2'd2)):(3'd5))}};
  localparam signed [4:0] p16 = {(~(3'd3)),(((2'd0)?(-2'sd1):(4'd8))^~((4'd14)!==(2'd2))),((5'd8)|(^(5'd24)))};
  localparam signed [5:0] p17 = (5'sd11);

  assign y0 = ((5'd15)!==({1{{1{(~&a2)}}}}>=$signed((~(4'd14)))));
  assign y1 = $unsigned(((((a3>>>b2)<=(p3^~p0))>>>((-b1)<$signed(b3)))<<<($signed((~^a5))%a4)));
  assign y2 = {(~&(!((a4<p9)=={p7})))};
  assign y3 = ({1{((a0?p6:p15)?(2'd3):(4'd6))}}<($signed((^{$unsigned(p5)}))));
  assign y4 = (-4'sd2);
  assign y5 = ((p9?p10:p2)?(-a4):(p1?p16:p0));
  assign y6 = (-2'sd0);
  assign y7 = $unsigned(((~|b1)&{p9,b0,a3}));
  assign y8 = ((-(($unsigned(b3)^$unsigned(a3))<(+$signed((b2+a5)))))|((-$unsigned((p5|a2)))>>$unsigned((~|(~|a4)))));
  assign y9 = (&(&(((b3|a0)!==(~^(~^a3)))^(-(!(3'd1))))));
  assign y10 = {{((p4<<<a2)?(a2?p4:b5):(4'd5))},(6'd2 * (b1<<p8))};
  assign y11 = (p7?a0:p4);
  assign y12 = (((b3?p7:a5)^(b4<<<b5))>>((b0+b5)?(b0&&a3):(|p0)));
  assign y13 = (~^(~|{((a5===a4)===(b3&&a1)),(~(-{p2,p8,b5}))}));
  assign y14 = {1{(5'd11)}};
  assign y15 = {(!{(!(~{(+a4),(a5?b2:b1)}))})};
  assign y16 = (((b1===b4)<<<(a3*b3))===(4'sd1));
  assign y17 = $signed($unsigned(($unsigned({4{b4}})<={4{b4}})));
endmodule
