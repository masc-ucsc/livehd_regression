module expression_00536(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(~^((2'd2)?(5'd15):(3'sd3)))},{((3'd4)>>>(4'sd1)),((5'sd9)||(5'd1))},(&((~(3'd3))<<((-2'sd0)?(3'd7):(2'd3))))};
  localparam [4:0] p1 = (-5'sd9);
  localparam [5:0] p2 = (((-3'sd1)*(3'sd2))<=(~(3'd0)));
  localparam signed [3:0] p3 = ((4'd12)?(~(3'd2)):{(-2'sd1),(3'sd0),(2'sd1)});
  localparam signed [4:0] p4 = {({(3'd7),(2'sd1),(-2'sd0)}>>(6'd2 * (5'd9))),{((4'd7)&(2'sd1)),((3'sd0)<<<(2'd1)),((-4'sd7)<=(-4'sd3))}};
  localparam signed [5:0] p5 = ((+(!((~^((-2'sd1)&(4'd2)))<<<((2'd3)<<<(-2'sd1)))))^~(~(~(~^{3{((5'd1)-(-2'sd0))}}))));
  localparam [3:0] p6 = {((5'sd7)^~(4'sd1)),((-5'sd6)>>(4'sd4)),((3'd3)^(4'd12))};
  localparam [4:0] p7 = (6'd2 * ((2'd1)<(3'd7)));
  localparam [5:0] p8 = ((((-4'sd2)&(-2'sd0))|((4'd9)>>>(3'd7)))||(((-3'sd3)===(5'd1))&&((5'd10)-(4'd6))));
  localparam signed [3:0] p9 = {3{{4{(4'd12)}}}};
  localparam signed [4:0] p10 = ((+(~|({3{(3'd1)}}^(5'sd4))))<=(2'sd0));
  localparam signed [5:0] p11 = ({{(-2'sd0),(5'sd13)}}|(~|{(5'd17),(3'd2)}));
  localparam [3:0] p12 = ((-2'sd1)?((2'd1)?(5'd10):(4'sd3)):((3'sd2)?(3'sd2):(2'sd1)));
  localparam [4:0] p13 = (((!(3'd0))*((4'd9)<=(5'sd1)))?((4'd2 * (5'd4))&&(~(2'd2))):(((3'sd1)<=(3'sd2))<<((3'd4)-(4'd5))));
  localparam [5:0] p14 = (5'd29);
  localparam signed [3:0] p15 = {{(4'sd5),(-5'sd7)},((4'd11)<(5'd21)),((4'sd4)^~(-4'sd4))};
  localparam signed [4:0] p16 = (5'sd7);
  localparam signed [5:0] p17 = (((-3'sd0)>>(5'd9))?((-5'sd2)?(4'd8):(5'd19)):((3'd1)?(4'd13):(-3'sd3)));

  assign y0 = (-2'sd0);
  assign y1 = {((p8<<a3)+{3{p17}}),((~|(b5|p14))-{a4,p2,p5})};
  assign y2 = {({{2{{4{(p4+b3)}}}}})};
  assign y3 = ({3{p9}}?(p4>p1):(p10?p5:p11));
  assign y4 = (((p15%p5)?(4'd3):(p9<p16))?((p4>a0)?(5'sd8):(4'sd0)):((3'sd3)));
  assign y5 = {4{{2{p1}}}};
  assign y6 = {(!$unsigned($signed((($unsigned($unsigned((|(|{(^(~{b5})),$unsigned((&(!b5))),{(b1),(&p11)}})))))))))};
  assign y7 = ((~&(~|{1{(b5^~b0)}}))!=((&(~a4))^{4{a0}}));
  assign y8 = (+(~&(^b1)));
  assign y9 = (-(&((2'd3)<<(~(2'd3)))));
  assign y10 = (^(+(((-p9)?(b5?b0:b2):{p9})?(!(~|(2'd0))):{(-3'sd0),(-4'sd4),{a0,a0}})));
  assign y11 = ((4'd2 * (+{1{a2}}))|{1{(+((b4==a4)-{2{p3}}))}});
  assign y12 = ((+({b5,a2}===(~(a0>>a2))))<<((b2>a2)+(a1&&p5)));
  assign y13 = {1{{2{({1{p10}}==(~&a3))}}}};
  assign y14 = ((-2'sd1)%b3);
  assign y15 = {{a3},(|p1),(p8<<a4)};
  assign y16 = {3{((b4^p4)>=(b2!==a4))}};
  assign y17 = {3{({1{a0}}||(a3|p13))}};
endmodule
