module expression_00324(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(2'd1));
  localparam [4:0] p1 = ((~&(((3'd4)?(3'sd1):(-5'sd4))!==((3'sd1)*(-2'sd1))))?(~(6'd2 * ((3'd7)>>(4'd8)))):(((3'sd0)>>(5'sd11))%(-4'sd4)));
  localparam [5:0] p2 = (!(((-4'sd0)?(-2'sd1):(5'd29))>>(&(3'd1))));
  localparam signed [3:0] p3 = {{(5'd8),(2'd1),(-3'sd2)}};
  localparam signed [4:0] p4 = (~(5'd22));
  localparam signed [5:0] p5 = {{3{(3'd4)}}};
  localparam [3:0] p6 = ((4'sd3)?(3'd4):(5'd31));
  localparam [4:0] p7 = {{4{(4'd1)}},(&(|(4'd13))),{3{(-3'sd3)}}};
  localparam [5:0] p8 = ((!(2'sd1))?((5'd29)||((-2'sd0)==(4'd12))):((-(2'd3))?((5'sd11)?(5'sd13):(4'd15)):(^(5'd30))));
  localparam signed [3:0] p9 = {3{((4'd0)^(4'd5))}};
  localparam signed [4:0] p10 = (!({{(-3'sd3),(5'sd0),(2'd0)},{3{(4'd12)}},((-2'sd1)>>>(3'd0))}<(((-5'sd13)^~(2'sd1))<(~|(3'd5)))));
  localparam signed [5:0] p11 = (((~((2'sd1)>>>(4'd12)))>((2'd2)<<<(-4'sd6)))^~(((-2'sd1)?(5'sd15):(4'd2))?(^(-4'sd0)):(3'sd3)));
  localparam [3:0] p12 = ((!(4'd13))?(+(5'd22)):{4{(3'd5)}});
  localparam [4:0] p13 = {1{{(3'sd1),(4'd5),(5'd9)}}};
  localparam [5:0] p14 = {1{(4'd2 * ((4'd3)!=(5'd15)))}};
  localparam signed [3:0] p15 = (+(((4'sd0)==(2'd0))||(|(5'd5))));
  localparam signed [4:0] p16 = ({3{(-5'sd0)}}<<<((2'sd1)>>>(5'd5)));
  localparam signed [5:0] p17 = {1{(((5'd28)?(3'd3):(3'd6))?((2'd1)?(-5'sd11):(4'd2)):{3{(4'sd1)}})}};

  assign y0 = (5'd2 * $unsigned((p17^p5)));
  assign y1 = {{{p15,b5},(p2<p16),(2'd3)}};
  assign y2 = (^(2'd1));
  assign y3 = (2'd3);
  assign y4 = (5'sd9);
  assign y5 = {(~{p5,a3,p16}),(b1!=p9)};
  assign y6 = ({3{{$signed((b3)),$signed({a1,a1})}}});
  assign y7 = $unsigned((~((3'd7)>=(2'sd0))));
  assign y8 = {2{(^a4)}};
  assign y9 = ((a0?a4:b0)===(b2<a5));
  assign y10 = (&(~&(5'sd8)));
  assign y11 = (((p11?p10:p0)?(p14?p10:p17):(5'd22))^((b5>>>a0)?$unsigned(b2):(~&p5)));
  assign y12 = $signed((((-4'sd7)==={4{a0}})+((3'd1)>=(p7|p8))));
  assign y13 = (b3-a5);
  assign y14 = ((-((p7==a4)|(+a1)))+$unsigned(({p4,b2}==(p10-p10))));
  assign y15 = {(3'd0)};
  assign y16 = {3{(a1?b1:b3)}};
  assign y17 = {{(&{({a5,b3}!==(!(b5<<b4))),{{{{(+a3),(a3+b1)}}}}})}};
endmodule
