module expression_00644(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd0)<=(3'sd2));
  localparam [4:0] p1 = (!({4{(4'd13)}}?((3'd3)|(5'sd1)):{(3'd4),(4'sd3),(3'd7)}));
  localparam [5:0] p2 = (~|{4{(~^(4'd2))}});
  localparam signed [3:0] p3 = (~(((3'd5)?(2'sd0):(-5'sd13))<<<((-3'sd1)?(5'sd12):(-4'sd0))));
  localparam signed [4:0] p4 = ((~&(((5'd16)<<<(2'd3))^((5'sd15)>=(3'd1))))==={1{(((3'd2)>>>(5'd21))^((5'd20)<=(3'd2)))}});
  localparam signed [5:0] p5 = ((-4'sd2)?(3'd7):(-3'sd2));
  localparam [3:0] p6 = (!(5'sd1));
  localparam [4:0] p7 = ({1{((3'sd2)?(4'd11):(2'd0))}}?((3'd1)?(5'd1):(2'd2)):(-5'sd11));
  localparam [5:0] p8 = ((2'd1)>>(2'sd1));
  localparam signed [3:0] p9 = (3'sd0);
  localparam signed [4:0] p10 = (6'd2 * (~^{3{(2'd0)}}));
  localparam signed [5:0] p11 = (((4'd9)>>(5'd15))?(3'd6):(-5'sd4));
  localparam [3:0] p12 = ((((3'sd0)||(2'sd0))||{(5'd0)})||(~|({(5'd0)}!==(-4'sd6))));
  localparam [4:0] p13 = {3{(4'd8)}};
  localparam [5:0] p14 = ((~|(4'd8))==((5'sd7)>(-3'sd0)));
  localparam signed [3:0] p15 = (-2'sd0);
  localparam signed [4:0] p16 = ({{(5'd18),(2'sd0),(-5'sd5)},{(-3'sd3),(2'd1),(3'd3)}}-{{(-5'sd7)},(-3'sd0)});
  localparam signed [5:0] p17 = {(4'd2),(3'sd3),(2'd2)};

  assign y0 = (|(-((~^((~^b2)?(b0-a3):(+p5)))>>((b5%b2)^~(a5<<<a4)))));
  assign y1 = (~({a3,p12}<<(!(^a0))));
  assign y2 = (|$signed((~|{2{b1}})));
  assign y3 = (p6+b5);
  assign y4 = (({4{a2}}?(p10<<b3):(b3===a5))<{(^{p15}),{{p6,p2}}});
  assign y5 = $signed(((-3'sd3)));
  assign y6 = {1{{2{{3{p9}}}}}};
  assign y7 = ({1{p8}}|(~&p10));
  assign y8 = (&(((|{1{(6'd2 * a1)}})|{4{b2}})-(-5'sd0)));
  assign y9 = (6'd2 * (b1&a1));
  assign y10 = $unsigned((((p12/p12)?(b1^p11):(p13+p7))<<<$unsigned(((b1===a0)&(p2<=p2)))));
  assign y11 = (|{{(b4!==a3)}});
  assign y12 = (a3<=p0);
  assign y13 = (~(p13&&p7));
  assign y14 = ((2'd2)<<<((~(5'sd1))>>>(+(a2&&a2))));
  assign y15 = ((($signed(b5)===(a4|b4))<((~&p2)<=(|a3)))>{(b3!=b4),(~^{b1,b2,b0}),(b1&a1)});
  assign y16 = ((-(-4'sd5))?((3'sd3)!=(a3>>>p11)):(5'd5));
  assign y17 = (({b4,a3,p16}^(~|p16))?((p4?p1:p8)>>>(p6&p14)):((p15?a1:p0)==(p14|b4)));
endmodule
