module expression_00535(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^((^(~(&{(5'd0),(-4'sd3),(5'd18)})))<{{1{(4'sd7)}},{(2'd0),(3'd4)},(+(5'd11))}));
  localparam [4:0] p1 = {1{((2'd2)|(-4'sd4))}};
  localparam [5:0] p2 = ((&(((3'd4)<<<(4'sd6))-(~|(2'd1))))||(((3'sd1)<(5'sd6))!=((-3'sd3)*(2'sd1))));
  localparam signed [3:0] p3 = {2{((2'd1)|(3'd5))}};
  localparam signed [4:0] p4 = (-3'sd2);
  localparam signed [5:0] p5 = (((3'd5)&(4'd2))&((3'sd2)&&(-3'sd0)));
  localparam [3:0] p6 = ((+(((5'd3)===(-2'sd1))!==(&(-2'sd1))))^~{4{(3'sd1)}});
  localparam [4:0] p7 = {4{(-5'sd7)}};
  localparam [5:0] p8 = ((2'd1)>(((5'd25)>(4'd4))?(2'sd0):((5'd4)&(5'd17))));
  localparam signed [3:0] p9 = (((4'd7)?(-3'sd2):(4'sd0))?(((3'd4)?(4'd14):(5'd23))||((5'd17)>=(2'd3))):({4{(2'd2)}}||{(-4'sd3)}));
  localparam signed [4:0] p10 = ({{2{(4'd3)}}}?{2{(3'd1)}}:{1{(-2'sd1)}});
  localparam signed [5:0] p11 = (4'd5);
  localparam [3:0] p12 = (|(~^(-3'sd2)));
  localparam [4:0] p13 = {{(-3'sd2),(4'd2),(2'd0)},{(3'sd2),(-2'sd0),(2'd2)}};
  localparam [5:0] p14 = (|(^(|((4'd4)>>{(4'sd7),(4'sd0),(3'd7)}))));
  localparam signed [3:0] p15 = {(4'd5),(4'sd5)};
  localparam signed [4:0] p16 = ((((5'sd11)||(3'd7))!={4{(5'sd5)}})?((-5'sd14)?(3'd3):(-4'sd4)):((2'd2)?(3'd6):(2'd2)));
  localparam signed [5:0] p17 = (((-2'sd1)?(2'd0):(4'd14))?((~^(-2'sd0))&&(-(3'd3))):((5'd17)?(-3'sd2):(3'sd3)));

  assign y0 = (((3'd7)!=(b3&b1))>={(3'd6),(4'sd2)});
  assign y1 = (5'd2 * a0);
  assign y2 = (^{3{(a4<p6)}});
  assign y3 = (~&(((b4?b0:a0)?(!(a3?b4:b0)):{{b3,a3}})!==((5'd2 * a2)?(~^{a3,a5}):(3'sd2))));
  assign y4 = (p17|p6);
  assign y5 = (p13||p1);
  assign y6 = ((-3'sd2)<((b0<<p3)%a4));
  assign y7 = (p13/b5);
  assign y8 = {1{$unsigned(($unsigned((-4'sd5))-$signed((5'd9))))}};
  assign y9 = (((p2<=p3)+(a5!==b5))<<<$signed({p16,p5,p4}));
  assign y10 = ((3'sd0)&((!(4'd10))&(4'd3)));
  assign y11 = (4'd4);
  assign y12 = (|{1{(-3'sd1)}});
  assign y13 = ((b3<=b3)?(b4+a3):(a2==a2));
  assign y14 = (((p5?p4:b0)?(p3<p2):(!{a2,p3}))!=((p11^b0)?(4'sd2):(b1?b2:p12)));
  assign y15 = ((~(p13?p8:p5))?(a5?p5:p16):(3'sd2));
  assign y16 = (4'd2 * a0);
  assign y17 = ((!(^(((~&a2)-(~^a1))!=((^b1)&(p4^~p12)))))!=(!((+{a5,a1,b4})||{(-b2),{b3}})));
endmodule
