module expression_00333(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{((4'd1)&(2'd2))}};
  localparam [4:0] p1 = (^(~^{{((~^(+(2'sd0)))||((|(2'sd0))?(~|(4'd12)):(~^(4'd10))))}}));
  localparam [5:0] p2 = {4{(~{(5'd31)})}};
  localparam signed [3:0] p3 = {1{(2'sd1)}};
  localparam signed [4:0] p4 = {1{(-{(|{2{((-5'sd6)?(5'd4):(4'd6))}}),{1{(!(~{3{(3'd1)}}))}}})}};
  localparam signed [5:0] p5 = (-(~|(-2'sd1)));
  localparam [3:0] p6 = ((~|(-3'sd0))<<({3{(3'd0)}}===((4'd2)<<<(5'd25))));
  localparam [4:0] p7 = (~&(|(~&(~|(-2'sd0)))));
  localparam [5:0] p8 = {2{{4{(4'd9)}}}};
  localparam signed [3:0] p9 = ((4'sd3)>>{3{(4'sd0)}});
  localparam signed [4:0] p10 = (4'd2 * (&(~(5'd7))));
  localparam signed [5:0] p11 = {3{({3{(3'd6)}}&(2'd3))}};
  localparam [3:0] p12 = (5'd16);
  localparam [4:0] p13 = (!(~(&(4'd1))));
  localparam [5:0] p14 = ((((5'sd7)|(5'sd6))^(~(4'sd1)))||(((3'd3)||(3'd7))||((3'd4)>=(-5'sd14))));
  localparam signed [3:0] p15 = (((~(4'sd6))==(~|(-2'sd1)))?(((5'sd13)!==(5'd23))>(+(4'sd1))):{3{(~|(-3'sd2))}});
  localparam signed [4:0] p16 = ({3{(-5'sd1)}}&&((2'd2)!==(2'sd1)));
  localparam signed [5:0] p17 = ((&(!(4'd1)))?{2{(-3'sd3)}}:(^((5'd20)-(2'sd1))));

  assign y0 = ($unsigned(((~&(a0===b1))!=(a3>>a1)))!==(^((a1*b1)<=(~&(3'd0)))));
  assign y1 = (+{(p9?p12:p6)});
  assign y2 = (5'd26);
  assign y3 = ({4{p15}}?(6'd2 * $unsigned((p7>>b5))):((a5===b2)?(-4'sd2):(p7+b1)));
  assign y4 = ((((b1>>a3)>>(b5!=b2))>>((a4>>>b5)||(b0==a4)))===((~^(a1>>>a4))<<<((6'd2 * b2)<(~|b3))));
  assign y5 = $unsigned({1{(|{(-{(p16||p10),{p5,p17},{(~|p14)}})})}});
  assign y6 = {(&{p14,p11,p3}),{(p15==p9)},(|{p4})};
  assign y7 = {(p4>p0)};
  assign y8 = (-((~(~^(+$unsigned(((^p10)|(~a1))))))-$unsigned(((&(~^b0))*$unsigned((^p12))))));
  assign y9 = (~|(-5'sd15));
  assign y10 = (((b1?b1:a1)?(b2?a2:b0):(p3?b2:b5))?{{b2,a3,p7},(b5?a1:b3)}:{($unsigned(a0)?$signed(a0):(b3))});
  assign y11 = ((~|p3)<={b3});
  assign y12 = ((5'd21)?(5'sd11):(&(5'd20)));
  assign y13 = ((p3^~b1)%b4);
  assign y14 = (~^{3{(~&a5)}});
  assign y15 = (~(+(-(+(|(((4'd1)<<(b5?a4:p17))+(3'd3)))))));
  assign y16 = {{1{{$signed((+{3{a4}}))}}},((-(b5>b5))<<<{{1{b3}}})};
  assign y17 = ((a1>=b3)===(b5===a1));
endmodule
