module expression_00583(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd2 * (2'd2))^{4{(4'd4)}});
  localparam [4:0] p1 = ({2{((5'd28)&&(3'd5))}}<((3'd2)>={3{(5'd13)}}));
  localparam [5:0] p2 = (~|((~^(^(3'd4)))===(6'd2 * (5'd2))));
  localparam signed [3:0] p3 = {1{(({(4'd3),(-2'sd0)}&&{2{(5'd3)}})|{4{(2'd1)}})}};
  localparam signed [4:0] p4 = (((3'sd0)<<(3'd4))?((3'd7)||(2'd1)):((3'sd2)?(5'd29):(-5'sd4)));
  localparam signed [5:0] p5 = (!({2{(!(3'd3))}}>{1{(!(~^{4{(4'd14)}}))}}));
  localparam [3:0] p6 = {(2'd3),((^(5'd22))===((2'd3)&&(4'sd0))),(3'd4)};
  localparam [4:0] p7 = {{1{{(4'd2 * (4'd0))}}},{(~&{4{(-4'sd0)}})}};
  localparam [5:0] p8 = {((4'sd6)>>>(2'd0))};
  localparam signed [3:0] p9 = ((4'sd5)?(3'sd2):(2'd1));
  localparam signed [4:0] p10 = {1{((5'd3)?(5'd15):(-5'sd4))}};
  localparam signed [5:0] p11 = ((2'd1)-{3{(2'sd0)}});
  localparam [3:0] p12 = (&(~^{{3{((5'd16)>>>(3'd3))}},({3{(2'd3)}}==(~(-5'sd7))),{2{{(-4'sd0),(4'd14)}}}}));
  localparam [4:0] p13 = {3{{3{(2'd0)}}}};
  localparam [5:0] p14 = {1{{2{(4'd8)}}}};
  localparam signed [3:0] p15 = ((((3'sd1)===(4'd10))!=((3'd7)-(2'sd0)))!==((6'd2 * (2'd1))?((3'sd3)>>(-4'sd0)):{(2'sd0)}));
  localparam signed [4:0] p16 = (({4{(2'sd0)}}!==((3'd7)!==(-5'sd10)))?(4'd2 * {4{(2'd3)}}):((5'd7)?(4'sd7):(2'sd1)));
  localparam signed [5:0] p17 = (2'd2);

  assign y0 = (~|({(b1==b2),$unsigned({a0}),((a5>a3))}<({a0,b3,a5}!=(!(|(b4>>>b4))))));
  assign y1 = ((+{{a2},(a3^~a5),(-4'sd1)})===(3'sd2));
  assign y2 = (^b5);
  assign y3 = (!(-4'sd2));
  assign y4 = {2{a3}};
  assign y5 = (-($unsigned(p6)?(a3):(~a5)));
  assign y6 = {(!p15),{p6,p0}};
  assign y7 = (((p16<p5)+(~(p13>b4)))?((a3^b4)!==(b4<=a3)):(-4'sd1));
  assign y8 = ((^(|b2))>{(5'sd5)});
  assign y9 = (2'sd0);
  assign y10 = ($signed($signed(((p14)<=$unsigned(p11))))>$unsigned((($unsigned(p11)>=(a3)))));
  assign y11 = (p4||p13);
  assign y12 = ((~&$signed(((^a1)<<(b3?b0:b4))))?((|(^p0))==(~&(a3>>>b3))):((a0?a0:b5)?(p13?p8:b0):(p11>>a5)));
  assign y13 = (|(3'd6));
  assign y14 = (~^(3'd4));
  assign y15 = (~((+p4)!=(-b2)));
  assign y16 = ((a4&a4)?(a2+p17):(-3'sd1));
  assign y17 = (((~|(p4>>p1))?(2'd0):(!{2{p1}}))>>>((2'sd0)<=((a3?b3:p10)?(-a4):(p6|a4))));
endmodule
