module expression_00387(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(~|(^(~|(~|({(-4'sd6),(-5'sd7),(4'sd1)}+(!(~|((-3'sd2)+(5'sd13))))))))));
  localparam [4:0] p1 = ((5'sd11)?((-2'sd0)?(2'd1):(4'd13)):((3'd4)>>(4'd11)));
  localparam [5:0] p2 = ((((2'sd1)!=(-2'sd1))&((2'sd1)/(-2'sd1)))>>>(((3'd6)<=(2'd2))<=((4'd11)||(-4'sd3))));
  localparam signed [3:0] p3 = (~((|(2'd1))?(|(4'd15)):((3'd3)?(4'd8):(5'd11))));
  localparam signed [4:0] p4 = ((-3'sd1)>>(-5'sd14));
  localparam signed [5:0] p5 = ((~&(5'sd0))?(-(5'sd8)):((4'd13)^(2'd2)));
  localparam [3:0] p6 = (-2'sd0);
  localparam [4:0] p7 = ((3'd5)?(5'd26):(-5'sd2));
  localparam [5:0] p8 = ((-(^{{(5'd3)}}))&&(&({(5'd26),(2'sd1),(5'd24)}!=(5'd2 * (3'd3)))));
  localparam signed [3:0] p9 = {3{((-5'sd1)^(5'd0))}};
  localparam signed [4:0] p10 = ({3{((3'd2)?(3'd5):(3'd5))}}?(~|((2'sd1)?(2'd1):(2'd1))):(!(((3'd0)?(5'sd13):(2'd0))<=(!(5'd31)))));
  localparam signed [5:0] p11 = (!{4{{4{(2'd0)}}}});
  localparam [3:0] p12 = ({(4'd13),(4'd7),(+(4'd7))}>>(3'sd3));
  localparam [4:0] p13 = (4'd5);
  localparam [5:0] p14 = (+((+(~((5'd27)?(5'd28):(2'sd0))))?(~|(^((3'd4)?(3'sd1):(3'sd1)))):(~|((2'sd1)?(-2'sd1):(4'd2)))));
  localparam signed [3:0] p15 = ((((-2'sd0)*(-5'sd5))&((5'd15)%(-5'sd2)))>>(((-2'sd0)!==(5'd23))>((5'd10)>=(5'sd15))));
  localparam signed [4:0] p16 = (((2'd0)&(-2'sd0))<=((3'd7)>>>(5'sd12)));
  localparam signed [5:0] p17 = ({(-(-5'sd15))}&&{2{(-4'sd2)}});

  assign y0 = (({3{b1}}?(a0?b0:b0):{a5,p12,a4})|({2{{b2,b2}}}^~{{3{b0}},(b3?a1:a3)}));
  assign y1 = $signed((2'd0));
  assign y2 = (((a1>>b5)<=(b3))|(($unsigned(a1)-(p0-a5))));
  assign y3 = (((b0?b2:b2)?(p1?b2:b2):(~&b1))?{1{(&{2{(b1==b4)}})}}:{1{(-4'sd6)}});
  assign y4 = (^(b5===b4));
  assign y5 = (p9^~p12);
  assign y6 = (2'd0);
  assign y7 = {1{(-(~^((3'd7)>(-5'sd11))))}};
  assign y8 = (-(2'd3));
  assign y9 = {(a1==b5),{4{b2}},(!{a0,a5})};
  assign y10 = {$signed(({(|((~(p17<<<p14))))}<(^{$unsigned(b4),(p14&&a5),(b0|p15)})))};
  assign y11 = (((b3^p11)!=(~(~&a3)))?((-(a3/b2))>=(a5!=a3)):(!((~|(a3?a5:b1))||(a1<a3))));
  assign y12 = (a0!==a4);
  assign y13 = {2{{2{a1}}}};
  assign y14 = ((-4'sd1)|(-5'sd4));
  assign y15 = {{$unsigned(((p12?p10:p14)?{p17}:$unsigned(p12))),({(a3?p2:b3),{p12,a3},(p2?p16:p11)}),{$unsigned({a2,p16}),{b0,p17,p8}}}};
  assign y16 = (+p16);
  assign y17 = (~|((b5*a0)<(3'd6)));
endmodule
