module expression_00044(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(4'd6)};
  localparam [4:0] p1 = (((2'sd1)?(2'd0):(3'd3))^~((4'd14)<=(-3'sd1)));
  localparam [5:0] p2 = (4'sd5);
  localparam signed [3:0] p3 = ((((4'd1)&&(3'sd0))?{4{(4'd3)}}:(+(4'sd4)))?(!(((2'd2)?(5'd19):(2'd1))>>{2{(5'd19)}})):({3{(3'd4)}}&&((2'd3)&(2'sd0))));
  localparam signed [4:0] p4 = {3{{4{(-2'sd0)}}}};
  localparam signed [5:0] p5 = ((~|(2'sd1))||(-(2'd3)));
  localparam [3:0] p6 = {((4'sd5)?(2'd0):(-2'sd1)),((2'd3)^~(3'd1))};
  localparam [4:0] p7 = (-2'sd0);
  localparam [5:0] p8 = ({3{((4'sd0)>>>(3'd3))}}>>>{4{(5'd27)}});
  localparam signed [3:0] p9 = (&(2'd0));
  localparam signed [4:0] p10 = ((3'd3)?{1{((3'sd1)?(-4'sd4):(4'd12))}}:(-2'sd0));
  localparam signed [5:0] p11 = (~{4{(3'd0)}});
  localparam [3:0] p12 = {{(3'sd1),(-3'sd1)},{(5'd18)},{(-4'sd4),(5'd3)}};
  localparam [4:0] p13 = {3{(((2'd3)<<<(5'sd0))<{3{(3'd3)}})}};
  localparam [5:0] p14 = (|((((3'sd3)==(4'd15))>((-2'sd0)>>>(5'sd5)))>>(^{(5'd9),(2'd3),(5'd10)})));
  localparam signed [3:0] p15 = (((2'sd0)!==(5'd5))?((2'd3)+(5'd24)):(+(4'd10)));
  localparam signed [4:0] p16 = (((-5'sd0)?(5'd30):(-4'sd1))?((-4'sd7)?(3'sd2):(5'd2)):((5'sd2)-(-5'sd13)));
  localparam signed [5:0] p17 = (~&(~(!(|((4'sd0)>>>((-5'sd8)===(5'd8)))))));

  assign y0 = $unsigned((2'sd1));
  assign y1 = ({p2,p3,p0}?{2{p2}}:(b2?p14:p9));
  assign y2 = $unsigned((-4'sd5));
  assign y3 = $unsigned(($unsigned($signed((5'd24)))?(5'd9):((p16-p1)&(b0===b0))));
  assign y4 = (((a1<=b1)?(a5>>>a3):(b4>>a2))||({2{b0}}+(b3<<<a3)));
  assign y5 = (&{1{(((b2||a1)<=(&a3))^{3{a0}})}});
  assign y6 = (((p6<a0)/a4)<((b0&p9)/b5));
  assign y7 = {{(5'd3),{(p14)}},(5'd27)};
  assign y8 = {{(^(|{p8,p17,b4})),((a2?p14:p4)-(~&p5)),({b4}!==(b5?a4:a1))}};
  assign y9 = ({p17,p4}^(!p15));
  assign y10 = ((~&(6'd2 * p7))<<<(b1?a4:p7));
  assign y11 = ((!((p11<<p8)/(1+p4)))^(((~b0)!==(b2<<b5))!=((2'sd0)?(-5'sd1):(&p0))));
  assign y12 = (5'd2 * (a1===a0));
  assign y13 = (~|(((a1?p4:b5)-((^b1)))&(|((p12?p0:b3)|(b0||p1)))));
  assign y14 = (p5?p8:b5);
  assign y15 = (!({(~^(~&(b3<b3))),(&{(a2?a5:a5)})}<<<(~&(+(-{(~&(+a3)),(+{p14,b4,p11})})))));
  assign y16 = {1{((!$signed({a1}))?$signed({a4,p16,p14}):(~&{a3,p0,b0}))}};
  assign y17 = {1{{1{b0}}}};
endmodule
