module expression_00203(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((6'd2 * ((5'd3)<=(2'd3)))<<<((((3'd4)==(2'sd0))>=((2'd1)*(4'd5)))>=(((2'd2)!=(-3'sd3))&&((4'd4)===(2'd2)))));
  localparam [4:0] p1 = (|(((-(~^(4'd2)))||(-((5'sd9)<<(2'd2))))>>(&(((-4'sd1)>=(5'sd13))>(|((4'sd7)+(5'd28)))))));
  localparam [5:0] p2 = (4'd0);
  localparam signed [3:0] p3 = ((+((5'sd2)!==(4'sd2)))<<{3{(4'd10)}});
  localparam signed [4:0] p4 = (-(~|(3'sd3)));
  localparam signed [5:0] p5 = ({2{((-3'sd1)|(2'd1))}}!={4{{3{(2'd0)}}}});
  localparam [3:0] p6 = (&(4'd11));
  localparam [4:0] p7 = {4{(4'd13)}};
  localparam [5:0] p8 = {(5'd31),(3'd0),(4'd2)};
  localparam signed [3:0] p9 = (~|((|(^{({2{(-5'sd12)}}||{4{(4'd1)}})}))^{{(3'sd0),(5'd10),(3'd2)},{((5'd25)===(2'sd1))}}));
  localparam signed [4:0] p10 = ((2'd2)?(2'd2):(3'd0));
  localparam signed [5:0] p11 = ({{(-3'sd0),(-4'sd3)},{(3'd7),(2'sd0)}}<=({(-2'sd0),(-5'sd15),(2'd1)}>=((3'd0)&&(4'd7))));
  localparam [3:0] p12 = {{3{(4'd8)}},(2'd1)};
  localparam [4:0] p13 = (-{(5'd9),(-5'sd6)});
  localparam [5:0] p14 = {{(-4'sd6),(5'sd10),(2'd2)},{1{((5'sd10)?(-2'sd1):(-5'sd12))}}};
  localparam signed [3:0] p15 = {4{((4'd12)<<(2'd2))}};
  localparam signed [4:0] p16 = ((2'd1)<<<(5'd2));
  localparam signed [5:0] p17 = (-5'sd11);

  assign y0 = ((&{2{(+(-b4))}})>>{4{(~a0)}});
  assign y1 = (~^(-3'sd0));
  assign y2 = (((-3'sd3)!==(4'd2 * b2))>>(~(-(-a3))));
  assign y3 = ((((6'd2 * b1)<<(b0==a5))>={4{b1}})<({(p17==a5),{3{b5}},(b2<a0)}^{{1{a1}},{2{a0}},{b1,p4,b2}}));
  assign y4 = ({4{(a3==b2)}}===({4{b3}}&&(!(a1>>>b3))));
  assign y5 = {{(({p4}^(p7==p13))>=((a2||a1)===(b5>>>b3)))},(({p5,p8}^~(p4&&p6))>>>((p7>>p0)!=(p12<p1)))};
  assign y6 = {{(4'd2 * (p1?p13:p1))},(((-5'sd6)|(3'd4))&((p2?p9:p10)>(p9<<b1)))};
  assign y7 = (|(p12?b3:b1));
  assign y8 = {b4};
  assign y9 = ({3{a2}}?{(a2?b2:b3)}:{a1,a5});
  assign y10 = ({{(~^{{3{p6}},(-p17),(~|b1)})}}>(({1{b3}}>(~|p7))+({1{a3}}-{a1,b3,p6})));
  assign y11 = {3{{4{p7}}}};
  assign y12 = ({4{a1}}^(2'sd0));
  assign y13 = ((b4?b1:a2)?(b2?a3:p9):(p6<p17));
  assign y14 = {({1{{({2{a2}}!==(a4<a0))}}}<<<{({3{p17}}!={1{p14}})})};
  assign y15 = (&((a2%p16)&&(!(a3!=a2))));
  assign y16 = ((((p0))&(a3&a1))<=(4'sd7));
  assign y17 = {1{(!({3{b0}}==(&p15)))}};
endmodule
