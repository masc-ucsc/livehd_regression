module expression_00408(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{{3{(((5'sd8)-(3'd7))<={1{(4'd11)}})}}}};
  localparam [4:0] p1 = {{1{(5'd9)}}};
  localparam [5:0] p2 = (~&{2{((4'd8)!=(-5'sd13))}});
  localparam signed [3:0] p3 = (|(((-3'sd0)?(-2'sd0):(5'd29))?(~|(4'd5)):(+(4'sd0))));
  localparam signed [4:0] p4 = ((~|((2'sd1)?(5'sd1):(-5'sd7)))===(|(~((-5'sd13)<=(-4'sd7)))));
  localparam signed [5:0] p5 = ((2'd2)?({4{(5'd20)}}>>{(2'sd1)}):{4{(4'sd0)}});
  localparam [3:0] p6 = ((-{2{((4'd7)===(5'sd6))}})!={1{{4{(2'd3)}}}});
  localparam [4:0] p7 = ({1{(5'sd9)}}&&((-4'sd6)<<(-4'sd6)));
  localparam [5:0] p8 = ((6'd2 * (3'd3))?(+((4'sd5)?(4'd7):(-3'sd0))):(5'd15));
  localparam signed [3:0] p9 = {{(-(5'sd6)),((4'd9)?(3'd7):(4'd0)),((2'd1)?(3'sd0):(-4'sd6))},{((4'sd4)?(-3'sd3):(-3'sd0)),{(2'sd1),(-2'sd0)}}};
  localparam signed [4:0] p10 = {{3{((3'd6)?(5'd6):(-3'sd0))}},{1{((-2'sd0)?(2'd2):(-2'sd0))}},((^(2'd3))||((4'd5)?(5'd25):(-4'sd6)))};
  localparam signed [5:0] p11 = (((-3'sd1)>>(-2'sd0))>>>((-2'sd1)?(5'sd11):(4'sd1)));
  localparam [3:0] p12 = (({(5'sd9),(5'sd2)}?{(-4'sd4),(3'd0),(5'd16)}:{(4'd15),(-5'sd2)})-{((!(5'sd15))?((3'd3)<<<(5'd9)):((3'sd2)?(5'sd3):(2'sd1)))});
  localparam [4:0] p13 = ((2'd0)?(3'd0):(-4'sd5));
  localparam [5:0] p14 = {{{1{{(-4'sd5)}}}},{(5'd1),(3'sd3),(3'd4)},{3{(3'd1)}}};
  localparam signed [3:0] p15 = (4'sd4);
  localparam signed [4:0] p16 = ((|((4'd11)>(4'd8)))^((3'sd0)?(-3'sd3):(2'd0)));
  localparam signed [5:0] p17 = (4'sd5);

  assign y0 = ((~^($unsigned(a4)*(a3!=b5))));
  assign y1 = (+((((-p5)^(p17>=p3))^(~&(!(b2>>>p7))))));
  assign y2 = ({1{{3{(^(b5?b2:a2))}}}}^(3'sd1));
  assign y3 = ((b3-b2)=={b3,p3});
  assign y4 = {1{((a0<<<b2)+(a2<<b5))}};
  assign y5 = {{a2},{1{a4}}};
  assign y6 = (~^(~&(~&(|(~(!(+(-(+(|(-(~|(^(!(!(&p9))))))))))))))));
  assign y7 = (2'd0);
  assign y8 = ((a5&&p7)^~(4'd7));
  assign y9 = ((4'd6)<{2{a1}});
  assign y10 = ((p17?a4:b0)*(b5*b0));
  assign y11 = {(3'd0),((b4<<b2)!==(b1<<<a3)),(~(!(a1<=p5)))};
  assign y12 = ((a1&p7)+(+{1{p6}}));
  assign y13 = {(3'd5),{(5'd24)}};
  assign y14 = {$signed((((p1-p9))^(b5?a5:p13))),((3'd7)&&{1{$signed(p6)}}),{4{$unsigned(p15)}}};
  assign y15 = (~&(&((|(a4))?(!(~^p4)):(^{b0}))));
  assign y16 = {p2,p1,p16};
  assign y17 = ({p6,b2,b5}?(~&(a3<p15)):((a0===a4)&(a2===b4)));
endmodule
