module expression_00074(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({3{(2'd2)}}<<<{3{(-4'sd0)}})+((~|(3'sd1))==((3'd1)|(4'd8))));
  localparam [4:0] p1 = (^(-(!(|(-(3'd1))))));
  localparam [5:0] p2 = (!({1{(5'sd6)}}>=(5'd2 * (!(|(4'd2))))));
  localparam signed [3:0] p3 = (+(!((&((-5'sd12)==(4'sd6)))^(~&(~((5'sd14)<<<(-2'sd0)))))));
  localparam signed [4:0] p4 = (((~|{(5'd29)})&((4'd14)|(4'd5)))^{{(~{{(2'sd1)},{(3'd6),(3'd7),(-2'sd0)}})}});
  localparam signed [5:0] p5 = (3'd5);
  localparam [3:0] p6 = ((-2'sd1)!==(-5'sd3));
  localparam [4:0] p7 = ((-5'sd2)===(4'd8));
  localparam [5:0] p8 = (((4'd1)?(5'd26):(3'd7))?((3'sd3)&&(4'd14)):((3'd7)^~(2'd2)));
  localparam signed [3:0] p9 = ((-2'sd0)<<(-2'sd1));
  localparam signed [4:0] p10 = (((-2'sd0)<<(3'd1))>=((5'sd7)||(-5'sd13)));
  localparam signed [5:0] p11 = {3{(4'd8)}};
  localparam [3:0] p12 = ((5'd10)-(5'd23));
  localparam [4:0] p13 = ((4'd2)<<<(5'sd7));
  localparam [5:0] p14 = (2'd0);
  localparam signed [3:0] p15 = (-(!(5'sd15)));
  localparam signed [4:0] p16 = {{((5'd25)>>(-2'sd1)),(|(3'sd0))},{((-2'sd0)===(-5'sd11)),(~(4'sd3))}};
  localparam signed [5:0] p17 = (~&((^((4'd9)<<<{(2'sd0),(-2'sd0)}))>=(3'd6)));

  assign y0 = {3{({b0,b4,a2}===(-4'sd7))}};
  assign y1 = (b5%a0);
  assign y2 = (a3?b2:p4);
  assign y3 = (a3?b0:b3);
  assign y4 = (~(((p15-b3)?{1{a3}}:(b3&p0))));
  assign y5 = ({p4,p5}?{a1,b2}:{(6'd2 * a1)});
  assign y6 = (!({4{p15}}&&{3{p2}}));
  assign y7 = (({1{{(a3>=b1)}}}===((a4&&a4)&(b5&b0)))>>>{4{(b3!=a0)}});
  assign y8 = (~(+$unsigned((-(-3'sd1)))));
  assign y9 = ((((a1===b0)!=(a4?b4:b1))-(b2?b5:b0))===({(a5>>>b0)}?(a3<<a3):(a1|a0)));
  assign y10 = ({(5'd8)}?(b4?p14:p15):(5'sd3));
  assign y11 = $signed((~^(|$unsigned(((p4?p12:p4)?$signed($signed({p8,p16})):{$signed(a1),(+p2)})))));
  assign y12 = ((6'd2 * (a1===a0))^((5'd2 * a2)-(b4>>>b2)));
  assign y13 = (4'sd6);
  assign y14 = (~^(!(^(|((~(p14?p2:p6))?(~(p1*p5)):(-(-p11)))))));
  assign y15 = (((p8&p11)-{p13,p9})<<((a2!==b2)<={1{{p14,p17,b4}}}));
  assign y16 = ((&((+(~(!(~|b4))))>>>(!$signed((p12/a5))))));
  assign y17 = ($signed(({4{b2}}?(a5!==b0):(b2|p8)))||((|({1{b0}}!={a1}))^$unsigned(((b2<=b4)&&(b2?a5:b5)))));
endmodule
