module expression_00252(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-4'sd1)>>(5'd0));
  localparam [4:0] p1 = (-5'sd11);
  localparam [5:0] p2 = ((((-2'sd0)!==(4'd12))!==((2'd1)>=(3'd4)))?((-3'sd1)?(2'd3):(4'd10)):((5'd29)?(5'd6):(5'd22)));
  localparam signed [3:0] p3 = {3{(4'd2 * ((2'd0)-(5'd20)))}};
  localparam signed [4:0] p4 = {4{{3{(-3'sd3)}}}};
  localparam signed [5:0] p5 = {{(5'd27),(-4'sd4),(2'd1)},(4'sd4)};
  localparam [3:0] p6 = {1{((2'sd1)?(5'sd4):(-3'sd1))}};
  localparam [4:0] p7 = {(((5'sd13)?(2'd3):(2'd3))&&((3'd2)?(2'sd0):(2'sd1))),((4'd12)?(4'sd1):(3'sd0))};
  localparam [5:0] p8 = (({(5'sd0),(2'd1),(2'sd0)}<={3{(5'd16)}})!={3{(-2'sd0)}});
  localparam signed [3:0] p9 = ({2{((3'd7)>=(5'sd1))}}>>{1{({3{(4'd12)}}^~{3{(5'sd14)}})}});
  localparam signed [4:0] p10 = (2'd2);
  localparam signed [5:0] p11 = {3{(~&(|(~&(4'd7))))}};
  localparam [3:0] p12 = {3{(-((-2'sd1)>(4'd1)))}};
  localparam [4:0] p13 = ((((2'd3)&(2'd1))*((2'd2)-(3'sd2)))<((+(~&(-4'sd7)))+(3'sd0)));
  localparam [5:0] p14 = {{3{(3'd6)}}};
  localparam signed [3:0] p15 = ((-5'sd9)?((4'sd3)?(3'sd1):(2'd1)):(5'd31));
  localparam signed [4:0] p16 = ({(4'd2),(3'sd1),(3'd1)}^~{{(2'd3),(2'd0)}});
  localparam signed [5:0] p17 = (((3'sd3)>>>(4'sd0))>=((-4'sd3)>=(-3'sd0)));

  assign y0 = (a1^a2);
  assign y1 = ((-4'sd0)<=(4'sd7));
  assign y2 = (5'd18);
  assign y3 = ({1{(5'sd15)}}<<<(((4'sd0)||(5'd11))^(-(b5||p17))));
  assign y4 = (6'd2 * {1{(p1>=p8)}});
  assign y5 = {{{(a0>=p7)}},{{p10},{p14}},{{{4{p6}}}}};
  assign y6 = (|{(-4'sd1),(5'sd0),(+p9)});
  assign y7 = (~^(-((&$unsigned($signed({2{(!b2)}})))!==({3{a2}}&&(+(+b5))))));
  assign y8 = (2'sd0);
  assign y9 = (({{p4}}^~(a5?b5:b4))?((a0===b5)?(~|p4):(^p8)):(|((p5>=p5)<<<(+{p16,p13}))));
  assign y10 = (~&((a0?a3:a4)?(-a0):(a2?b3:a0)));
  assign y11 = {4{(((4'd2 * p14)!=(b0!=p17)))}};
  assign y12 = ((-4'sd4)^(a3>>>b4));
  assign y13 = {4{((b4&&a4)||$unsigned(a4))}};
  assign y14 = ((p17?p16:p12)>$unsigned(p1));
  assign y15 = (5'sd7);
  assign y16 = ((((p0*p17)^(p15!=p13))||((b2<<b1)===(a1&&b1)))>=(((p7^p8)*(p17!=p15))!=((p9^p1)%p7)));
  assign y17 = ((p9&&p6)*(2'd2));
endmodule
