module expression_00863(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd2 * ((5'd28)^~(5'd30)))-{3{((3'sd0)^(2'd1))}});
  localparam [4:0] p1 = {{((4'sd3)-(3'sd0)),((5'd1)&(-4'sd6))},{((3'd6)!=(4'd0))},((-(-3'sd3))-{(2'd3)})};
  localparam [5:0] p2 = (!{(~&{{(3'd6)},{(4'd10)},{(5'd28),(-4'sd6)}})});
  localparam signed [3:0] p3 = {({(2'd1),(-3'sd2),(4'sd5)}===((-2'sd1)<<<(4'sd0))),(&{(^(3'sd1)),{(5'd20),(5'd18)}}),(&(~(&(~|(-2'sd1)))))};
  localparam signed [4:0] p4 = ((5'sd13)<<(2'sd1));
  localparam signed [5:0] p5 = ({{((5'd20)<<(4'sd7)),((4'd6)==(4'd2))}}!==({2{(3'd5)}}-(4'd14)));
  localparam [3:0] p6 = ((~{1{(3'd2)}})&(5'sd2));
  localparam [4:0] p7 = {3{((4'd2)?(5'd12):(-4'sd1))}};
  localparam [5:0] p8 = ((((2'd3)!=(2'd0))||((-4'sd0)!==(-5'sd5)))-(((5'sd2)<=(2'sd1))/(-3'sd0)));
  localparam signed [3:0] p9 = (((4'd0)<<<(-2'sd0))>>{(2'd2),(-4'sd2)});
  localparam signed [4:0] p10 = (&((!((|(5'd13))<=((3'd2)^~(4'd11))))?({(4'sd7)}?((4'sd6)?(4'sd5):(5'd0)):(-3'sd2)):(+((-3'sd2)?(2'd2):(4'd11)))));
  localparam signed [5:0] p11 = ((-5'sd4)?((2'd1)^~(5'd0)):((3'd2)?(-2'sd0):(4'd8)));
  localparam [3:0] p12 = ({{(3'sd0),(5'd8),(3'd7)},{(5'sd15)}}<(+(!((-4'sd2)^~(3'd7)))));
  localparam [4:0] p13 = {2{((3'd1)^~(-5'sd6))}};
  localparam [5:0] p14 = ({2{{1{(4'd13)}}}}^~(((-4'sd0)!==(-2'sd1))!=(^(2'd0))));
  localparam signed [3:0] p15 = (3'd7);
  localparam signed [4:0] p16 = ((((2'd3)<<<(2'sd1))>=((-4'sd1)&(3'd4)))!=={2{{1{((-2'sd1)<=(4'sd4))}}}});
  localparam signed [5:0] p17 = {3{{{2{((2'd3)?(3'd3):(2'd3))}}}}};

  assign y0 = ({(a5)}!=(~&(b3-b4)));
  assign y1 = (~&((-4'sd7)?((b5?b1:a2)&(a5?b5:p17)):(|(&{b0,a0,b3}))));
  assign y2 = $signed($signed((b0&b2)));
  assign y3 = ({2{(p9||b3)}}>((p3?p5:p6)?(p2?p7:p3):(a3<<<p0)));
  assign y4 = $unsigned(($signed({(a5>b4),((a4||a3))})===((b5>>a3)&(b1|a5))));
  assign y5 = (^(~(+(^(p12>=b4)))));
  assign y6 = {4{((b2>a2)^(5'd2))}};
  assign y7 = ((((b2^~a1))>>$unsigned((p5?p14:a4)))&&((b1?p15:p9)>>>{p12,p12,p10}));
  assign y8 = ((((a4?p8:p11)<=(-2'sd0))?((a3|p5)*$signed(p17)):((a5?b1:p9)*(p7/b0))));
  assign y9 = (((b1?p6:p7)?{p13,b2,a3}:(5'd2 * p8))>>>(4'd5));
  assign y10 = $signed(($unsigned((5'd2 * (3'd5)))>>$unsigned((4'd12))));
  assign y11 = ((~|(b3^~p14))%p1);
  assign y12 = ({p8,a2,a5}?(b4?p6:p14):(p12?a0:p13));
  assign y13 = ($signed((((a0!==a1)<(a5*a0))===($signed((a5>=a4))))));
  assign y14 = ((-4'sd5)!=={(5'd28),$signed({a2,a3}),(b3!==a4)});
  assign y15 = (~&{1{{(~^p9),{3{a5}},(-b0)}}});
  assign y16 = (~|(^{3{(&(|{4{a5}}))}}));
  assign y17 = {({{a3,p6,a1}})};
endmodule
