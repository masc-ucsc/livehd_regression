module expression_00315(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd13);
  localparam [4:0] p1 = {4{(-2'sd1)}};
  localparam [5:0] p2 = ({(-(5'd12)),(!(5'd6))}|((-4'sd5)+((5'd21)>>(4'd7))));
  localparam signed [3:0] p3 = (4'd1);
  localparam signed [4:0] p4 = (((5'd2 * (5'd30))===((-5'sd15)!=(4'd12)))+(((5'd16)<(5'sd3))/(4'sd5)));
  localparam signed [5:0] p5 = (!(&(~(3'sd2))));
  localparam [3:0] p6 = {(!{1{{(3'd3),(4'sd6),(-3'sd1)}}}),{1{(~^(+(-4'sd4)))}}};
  localparam [4:0] p7 = ((4'sd4)<=((-4'sd1)<<(2'd1)));
  localparam [5:0] p8 = ((-3'sd3)&(3'd6));
  localparam signed [3:0] p9 = ((-5'sd7)?(4'd6):(4'd11));
  localparam signed [4:0] p10 = (~|(((-3'sd2)?(2'd1):(2'sd1))-(-2'sd1)));
  localparam signed [5:0] p11 = (((2'd3)<=(2'sd0))?((3'd1)<<(-4'sd5)):((4'sd3)>=(-4'sd2)));
  localparam [3:0] p12 = (4'sd1);
  localparam [4:0] p13 = (3'd4);
  localparam [5:0] p14 = {{(|(4'd2)),{(4'sd3)},{(5'sd14)}}};
  localparam signed [3:0] p15 = ((4'd14)<(-4'sd6));
  localparam signed [4:0] p16 = ((5'sd1)^(4'd9));
  localparam signed [5:0] p17 = {3{(4'd5)}};

  assign y0 = (((4'sd7)^(p17|p8))?{1{(5'd5)}}:{(~&p6),{3{p9}}});
  assign y1 = {(-5'sd2),{p5,p10,p6}};
  assign y2 = (4'd14);
  assign y3 = {1{{{1{$unsigned({$unsigned($signed({p16,b2,b2}))})}},{4{(a0?p9:a1)}},{{{p10},{b2},{b0,p9}}}}}};
  assign y4 = (~&((p10>>p4)?(+(!p16)):(p0&&p10)));
  assign y5 = {((b3-a2)==(b5!==b5)),((|b5)&$signed(a1)),{2{{4{b0}}}}};
  assign y6 = (((b0||a5)?(2'd2):(~^a0))===(&{4{b4}}));
  assign y7 = (&(~|(!(&(~|((!(~^p0))/p12))))));
  assign y8 = (^(-5'sd6));
  assign y9 = (~^(^{4{{2{(-b1)}}}}));
  assign y10 = (|(p16?p11:p12));
  assign y11 = (5'sd4);
  assign y12 = {((a0<<b4)?(b5^b5):(b1||a5)),(2'd0)};
  assign y13 = ((($unsigned(a5)==={a5,b3,a4}))?((b1?a1:b1)>>>(b1<<p7)):{(p13?b5:p14),{p4,p2},$signed(b2)});
  assign y14 = ({(p6<p2),{p7,p3},(p1!=p16)}!={(p11<p11),(b1>=p4)});
  assign y15 = (5'sd11);
  assign y16 = ((b5?b2:a2)?(b5>b5):(b5!=a4));
  assign y17 = (((~|(p14?a0:a1))||((a1>b5)!==(b4|a5)))+{2{(~^{4{p1}})}});
endmodule
