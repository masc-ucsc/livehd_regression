module expression_00274(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd11)?(-4'sd4):(-5'sd7));
  localparam [4:0] p1 = (4'd1);
  localparam [5:0] p2 = (((4'd6)||(5'd16))?((2'd2)?(2'sd0):(5'd12)):((3'd6)?(4'sd0):(4'sd5)));
  localparam signed [3:0] p3 = (((+(-4'sd5))<=(+(-5'sd3)))<=(((-4'sd2)?(5'd20):(4'sd1))?((4'd3)||(-2'sd0)):(5'd12)));
  localparam signed [4:0] p4 = (3'd7);
  localparam signed [5:0] p5 = ((~^{2{(+(2'd2))}})<<<(+{{1{{(5'd20)}}}}));
  localparam [3:0] p6 = ((-4'sd6)?(2'd1):(2'd1));
  localparam [4:0] p7 = (4'sd3);
  localparam [5:0] p8 = {({(-4'sd1),(3'd4)}?{2{(-2'sd1)}}:((3'sd0)?(4'sd6):(2'sd1))),{((3'd3)?(-5'sd11):(3'd6))}};
  localparam signed [3:0] p9 = (((-4'sd1)>(5'sd8))===((2'd2)==(2'd3)));
  localparam signed [4:0] p10 = (4'd13);
  localparam signed [5:0] p11 = (((2'd2)<<(-4'sd3))<(2'd3));
  localparam [3:0] p12 = (3'd3);
  localparam [4:0] p13 = {4{((2'd0)?(-3'sd2):(-5'sd4))}};
  localparam [5:0] p14 = ({{1{(-2'sd1)}},{(3'd0),(5'd4),(5'd16)}}+({(2'd1),(2'd2)}>>((3'sd1)&(-4'sd5))));
  localparam signed [3:0] p15 = {{(3'sd2),((4'd9)^~(5'd10))},(~&(3'd0)),({(3'd7),(3'sd0)}?{(-5'sd1)}:{1{(-3'sd0)}})};
  localparam signed [4:0] p16 = {1{(|((~&{4{(4'sd0)}})==(|({2{(-5'sd14)}}^~{3{(4'sd7)}}))))}};
  localparam signed [5:0] p17 = (5'd2 * (4'd13));

  assign y0 = (~$signed(((((-$unsigned((~|a4)))+(~|(&(p1>>p8))))))));
  assign y1 = ((|(-p17))?((^a3)):(p5?b0:p13));
  assign y2 = (&{b2,a3,b3});
  assign y3 = ((-((b5?b3:a5)===(a3^~b2)))?(|{3{b0}}):(~^((p7?a4:a4)>>(b4&&p6))));
  assign y4 = ($signed(b2)?{p11,a5,p12}:$unsigned(b0));
  assign y5 = {3{{a5,p16,p14}}};
  assign y6 = {$unsigned($unsigned({{b0,p10,p16}})),$signed(($signed((p9))&&(p3|p10))),((a0!==b5)>$unsigned((a3|p2)))};
  assign y7 = {4{p2}};
  assign y8 = ((p15>>>p7)<<<{1{{p9,p10,p3}}});
  assign y9 = (5'sd10);
  assign y10 = (($unsigned($unsigned((p11<<<p15)))<<(^(~&(p4^~p11))))<=((a3&p15)?$unsigned($unsigned(p10)):(&(p16))));
  assign y11 = (~^p8);
  assign y12 = {(4'sd2),(({2{b3}})!=((b1===a4)==={3{b1}}))};
  assign y13 = (|(-(~&(^(&(~^(&(-(~|(-(-(~|p5))))))))))));
  assign y14 = (~|{(&(p15>p4)),(a5^b3),(b5?p1:p7)});
  assign y15 = ($signed((p15&a4))?((b0?b2:p9)<<(b2===b0)):(|(p11>>>p3)));
  assign y16 = (((3'd4))?(-3'sd0):(5'd14));
  assign y17 = (((a5+b3)!=={a3,a1})^({a0,a4}?(4'd6):(3'sd2)));
endmodule
