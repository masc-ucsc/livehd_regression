module expression_00038(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~(~|(3'sd3)))!=(~|(&(5'd16))));
  localparam [4:0] p1 = (-4'sd4);
  localparam [5:0] p2 = (|(~&(!((3'd4)^~((-5'sd2)&(2'sd1))))));
  localparam signed [3:0] p3 = (((-2'sd1)-((-5'sd10)?(5'd23):(4'sd6)))?(~|((5'sd14)<(-2'sd1))):{1{(~|(~|(2'd1)))}});
  localparam signed [4:0] p4 = ({1{{4{(3'sd2)}}}}?((4'sd7)?(4'd5):(4'd9)):((-4'sd0)>>(2'sd0)));
  localparam signed [5:0] p5 = ({2{(4'sd0)}}?({4{(-5'sd12)}}<<<((-2'sd1)<<(2'd3))):(-5'sd14));
  localparam [3:0] p6 = (~(-3'sd3));
  localparam [4:0] p7 = (!(3'sd0));
  localparam [5:0] p8 = (3'd6);
  localparam signed [3:0] p9 = {(+{3{(5'd2 * (5'd12))}})};
  localparam signed [4:0] p10 = {3{{1{((3'd6)?(5'd18):(3'sd0))}}}};
  localparam signed [5:0] p11 = ({2{((4'd13)<<(5'd7))}}^(&{(4'd2 * (2'd0)),{3{(5'd15)}}}));
  localparam [3:0] p12 = ((~(2'd1))<<((2'sd0)&(3'sd1)));
  localparam [4:0] p13 = (^(~(((-5'sd8)===(-2'sd1))%(3'd0))));
  localparam [5:0] p14 = (-({(5'd20),(-2'sd0)}>>{(4'd4),(4'd13)}));
  localparam signed [3:0] p15 = {(((-3'sd1)?(5'd1):(-4'sd5))?(5'd2 * (2'd3)):((-5'sd10)?(4'd2):(3'd1))),(5'd2 * {(2'd2),(2'd3)}),(((-3'sd3)>>(4'sd7))+((-2'sd1)>>>(-3'sd1)))};
  localparam signed [4:0] p16 = {2{(((2'sd0)>>(-5'sd2))|((3'd0)<(5'd15)))}};
  localparam signed [5:0] p17 = ((-2'sd1)&(^(-(5'd30))));

  assign y0 = {2{({2{{4{p6}}}})}};
  assign y1 = (3'd7);
  assign y2 = ($unsigned((~^(((p13==a1)>=(p2>>b0)))))^(~|((5'd2 * p6)|(p12^p6))));
  assign y3 = (((^b5)<(a1?a4:b5))?((+a0)<<(b3?p12:b2)):((p16?a1:p12)<<<(!a2)));
  assign y4 = ((-(+(!(a5<=b4))))<<((-4'sd2)^(b4&&a2)));
  assign y5 = {(({a1,a2,b3}>>>(4'd15))<={(p13+b1),(a3<<p8)})};
  assign y6 = (p2?p9:p4);
  assign y7 = (((-b2))|(b1?a4:b3));
  assign y8 = (((b3?a4:a0)?{3{a2}}:(a5?p6:b1))?(3'd7):((5'sd8)?{2{p8}}:(-2'sd1)));
  assign y9 = (4'd3);
  assign y10 = (+((-(&(~|((a1<<b3)==(~^a2)))))<(((a2&&b2)==(a4>=a2))&&((p7<p15)^(!b4)))));
  assign y11 = (~^(((~|p5)%p11)<<<(^(~^(~|b4)))));
  assign y12 = $signed((4'd3));
  assign y13 = (|(^(~|(2'sd1))));
  assign y14 = (~^$signed(((|(5'd9))/b4)));
  assign y15 = (p5>>b2);
  assign y16 = (((p11<=a4)?(~(^p10)):(p13?a4:p17))>{2{{{4{p6}},(b1-p8)}}});
  assign y17 = (((^$signed($signed((~|(~($unsigned(a2)<=(a4)))))))||(-(~$signed(((~^(~^a2))|$signed((b1^b3))))))));
endmodule
