module expression_00563(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{({2{(~^(2'sd0))}}-(~|(4'd6)))}};
  localparam [4:0] p1 = {(~(-4'sd5)),(3'd5)};
  localparam [5:0] p2 = (&(~(^({(-4'sd0)}!=((4'sd2)^~(4'sd2))))));
  localparam signed [3:0] p3 = (({(2'sd0),(-3'sd1)}<((4'sd0)&(4'd10)))?{((4'd11)>>>(4'd8))}:(6'd2 * ((4'd10)?(5'd0):(4'd11))));
  localparam signed [4:0] p4 = {(-{4{(!(5'd4))}})};
  localparam signed [5:0] p5 = {({3{(4'd0)}}?{(2'd3),(4'sd2)}:{(4'sd3),(5'd19),(2'd1)}),(|((5'd15)?(4'd12):(2'd1)))};
  localparam [3:0] p6 = (((4'd10)<(2'd2))-(^(5'd7)));
  localparam [4:0] p7 = (((~&(2'd3))!=((2'd2)>>>(-3'sd0)))!==(((3'd5)==(3'd1))>((-5'sd12)?(4'd7):(3'sd3))));
  localparam [5:0] p8 = ((3'd1)>(-2'sd1));
  localparam signed [3:0] p9 = (3'd3);
  localparam signed [4:0] p10 = {{(5'd2 * (4'd6)),{(-2'sd1),(4'sd7)}},(((-4'sd1)<=(3'd0))&((4'd3)>=(4'd9))),(((4'd14)<=(3'sd3))|((3'd3)>>(-3'sd3)))};
  localparam signed [5:0] p11 = ({4{(-5'sd11)}}^~(&(~&((-5'sd9)^(3'd1)))));
  localparam [3:0] p12 = ((3'd6)!==(2'd0));
  localparam [4:0] p13 = ((-(((-2'sd1)>>(3'd7))^~((3'd0)!=(2'd0))))>=(((2'd0)!==(4'd15))*((-4'sd7)?(2'd2):(2'sd1))));
  localparam [5:0] p14 = (((-2'sd0)&&(4'd9))<<((3'sd2)<(4'd4)));
  localparam signed [3:0] p15 = {{{{(2'd2)},(5'd6)}}};
  localparam signed [4:0] p16 = (~&({{(4'd8),(-3'sd3)},((3'd2)!=(-2'sd0)),((4'd10)?(3'sd0):(-5'sd1))}<<<({(4'sd5),(-4'sd0),(5'sd6)}!=((5'd12)!=(2'd1)))));
  localparam signed [5:0] p17 = ({1{(^{1{(4'd3)}})}}<<{3{(4'd13)}});

  assign y0 = (-4'sd2);
  assign y1 = {4{(|p3)}};
  assign y2 = (~|(&(({a2,b2}?(5'sd15):(b2?b4:p0))+((b5?b1:b2)<(a4|b0)))));
  assign y3 = {1{(5'sd14)}};
  assign y4 = (-((p6^~p15)));
  assign y5 = (~((~&(b1?b2:a5))?{{p6,b4},{4{p13}},(~|p0)}:(+{{1{(p4?p9:p15)}}})));
  assign y6 = ((p11^p17)*(b5===a0));
  assign y7 = {((p12<<<p13)!=(|a0)),((a2<b2)!==$unsigned(b1)),{({p13}&{p4,a5,p5})}};
  assign y8 = {{({{b5,b1,a1}}>>(~^{b1,b0})),{{b1,b5,a0},(b2^~b5),(p9<<b0)},({(b1|p10)}-(a4>>>a4))}};
  assign y9 = {(~(!$unsigned((a2^b3)))),$unsigned({(&a0),{b2},{b2}}),(-$unsigned((~^(~(b0^~a5)))))};
  assign y10 = {3{{4{(p8?b3:b5)}}}};
  assign y11 = {p10,b4};
  assign y12 = ({1{((p6<<<b0)?(~^{a2,p9}):{2{p10}})}}&{({4{a1}}?(-(a0?p11:b2)):(p12?p1:p16))});
  assign y13 = (-5'sd8);
  assign y14 = (2'sd1);
  assign y15 = (+{((a0?a2:a1)<<<(~^(a0?a5:a2))),(&(&((+b4)?(~b1):(b1!=a0))))});
  assign y16 = (+(-(^(|((p10?p13:p6)?(|p11):(~&p1))))));
  assign y17 = ((2'sd0)+(5'd24));
endmodule
