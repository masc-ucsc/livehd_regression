module expression_00875(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd2 * ((3'd5)==(2'd0)));
  localparam [4:0] p1 = ((5'd26)?(4'sd5):(2'sd1));
  localparam [5:0] p2 = (5'sd2);
  localparam signed [3:0] p3 = (((3'd2)<<(4'd0))?{(4'd6),(3'd7)}:{(-5'sd11),(-5'sd7)});
  localparam signed [4:0] p4 = {(4'sd0),(5'd13),(2'd1)};
  localparam signed [5:0] p5 = {((5'd2 * ((4'd9)^(4'd3)))==={{((4'd7)<<<(4'sd2)),{(4'd5),(-4'sd0)},{(2'd1),(5'd27),(3'd1)}}})};
  localparam [3:0] p6 = (^(+(&(~^(+(-(!(~&(~|(~&(-(~^(-(~&(~(3'sd3))))))))))))))));
  localparam [4:0] p7 = ({(5'd22),(-4'sd3),(2'd0)}?(~^(5'd24)):(~|(5'd28)));
  localparam [5:0] p8 = (~&(-5'sd6));
  localparam signed [3:0] p9 = ((((4'd11)==(5'd20))<<((2'd3)<=(3'sd2)))^{{(~^(4'sd7)),(~(-2'sd0)),{1{(5'd3)}}}});
  localparam signed [4:0] p10 = (6'd2 * {3{(5'd17)}});
  localparam signed [5:0] p11 = ((4'd3)&&(~&(3'sd3)));
  localparam [3:0] p12 = (((4'sd1)==(5'sd10))+{4{(3'sd1)}});
  localparam [4:0] p13 = (3'd0);
  localparam [5:0] p14 = ({(2'd3),(5'sd3),(5'sd12)}?((-5'sd13)>>>(2'sd1)):((2'sd0)?(5'd1):(2'sd1)));
  localparam signed [3:0] p15 = ((-(-5'sd6))?{2{(4'd1)}}:(~(4'd3)));
  localparam signed [4:0] p16 = ((4'd8)===(4'd7));
  localparam signed [5:0] p17 = (3'd2);

  assign y0 = {1{(5'd16)}};
  assign y1 = {(p2==p15)};
  assign y2 = (-((((a5?a2:b4)-(a0>>b1))===(-3'sd1))));
  assign y3 = ((p3?b1:b3)&(b4?b4:a2));
  assign y4 = (5'd31);
  assign y5 = ({1{(|a1)}}<(~^(a3?b5:a0)));
  assign y6 = (((~(~|b3))!==(6'd2 * b0))^({2{a0}}===(~&(~|b3))));
  assign y7 = ({({b4,p12,a5}<=(2'd0))}>=((a3^p8)|(4'd12)));
  assign y8 = (((a4?b3:p11)?(+(p2?b0:a5)):(^(b4!=b1)))!=$signed($unsigned(((a4?b4:b0)!==(&(a4?a2:a5))))));
  assign y9 = (p15||a3);
  assign y10 = {(2'd0),(4'd7),(+((p7^a2)+(b5>a3)))};
  assign y11 = (4'd2);
  assign y12 = (~&((5'd21)));
  assign y13 = ((p13^p16)-{p1,p12});
  assign y14 = {2{{2{{p3,b0,b1}}}}};
  assign y15 = {4{p4}};
  assign y16 = (b1>>a1);
  assign y17 = {((a4?a0:p12)-(b0?b0:p17)),{(b1-b1),(p9<p15)},((a3>>>a2)!==(a2?b0:b2))};
endmodule
