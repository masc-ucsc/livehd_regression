module expression_00608(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-4'sd5)?(4'd15):(5'd13))!=={(-3'sd1),(4'sd2)})>=(4'd1));
  localparam [4:0] p1 = (&(~|{(~((5'sd6)>>>(-5'sd3))),(((5'sd12)?(2'sd1):(3'sd3))>=((4'd13)+(4'd10))),{(2'd2),(2'd2),(5'd31)}}));
  localparam [5:0] p2 = (((-5'sd9)+(5'd0))<<<((2'sd1)?(-5'sd8):(5'd26)));
  localparam signed [3:0] p3 = {1{((5'sd13)&((3'd1)&&(4'd7)))}};
  localparam signed [4:0] p4 = (((4'sd4)>=(4'sd2))<(4'd9));
  localparam signed [5:0] p5 = ((~&((3'd0)?(-5'sd10):(4'sd6)))?(|(4'd12)):{1{(~|(4'd3))}});
  localparam [3:0] p6 = {4{{{(2'd2),(3'sd3),(5'sd9)},{1{(2'd3)}}}}};
  localparam [4:0] p7 = ((-2'sd0)?(2'sd0):(5'd17));
  localparam [5:0] p8 = {{1{{3{((-2'sd1)<(3'd6))}}}},{{(4'd0),(2'd1),(3'd5)},(-(4'd6)),(!(4'd9))}};
  localparam signed [3:0] p9 = (-((5'd10)>>>(3'd5)));
  localparam signed [4:0] p10 = (((|(3'sd1))>>>((3'd5)<<<(-4'sd3)))===(5'd2 * ((5'd31)&(5'd10))));
  localparam signed [5:0] p11 = {1{{1{{{{((2'sd0)?(4'd9):(-5'sd7)),{(3'sd2),(3'd3)}}}}}}}};
  localparam [3:0] p12 = ((((2'd0)|(4'd6))==(3'sd2))<=((-5'sd12)===(2'd1)));
  localparam [4:0] p13 = ((^(3'd5))==={1{(3'd2)}});
  localparam [5:0] p14 = ((3'd1)?{(5'd21),(-4'sd7),(5'd30)}:{(4'd4)});
  localparam signed [3:0] p15 = ((((4'sd0)<<<(-4'sd4))^~((2'd3)>=(-5'sd7)))&({2{(4'sd4)}}&(4'd2 * (3'd3))));
  localparam signed [4:0] p16 = ((4'd2 * (5'd22))>={4{(2'sd1)}});
  localparam signed [5:0] p17 = (~^{(~|(~&((2'd0)===(4'd2)))),((-(3'd0))+((-2'sd0)>>>(-3'sd2)))});

  assign y0 = (({{1{b5}},(p12?a2:p14)}<=((b3?a1:b2)||{a0,b1}))^~{(p15?b4:b1),(b1<<b4),(b3&p9)});
  assign y1 = ({(p1!=p12),{p11}}?(&{3{p16}}):($unsigned((p4|p0))));
  assign y2 = (^(3'sd2));
  assign y3 = ((^({1{(b5^p11)}}^(!(p5^b0)))));
  assign y4 = (a0?p4:p12);
  assign y5 = {3{{4{{3{b0}}}}}};
  assign y6 = $unsigned((((p0+p13))));
  assign y7 = (4'd10);
  assign y8 = (3'd5);
  assign y9 = (3'sd2);
  assign y10 = {b1,p2,p9};
  assign y11 = (~|$signed(((|(p13<=p12)))));
  assign y12 = {((a2>>>p6)),(a3^p13),((p6))};
  assign y13 = (|(((!{a4})<<<{b3,a0,a5})<={{(p10?b5:a0)},(b0?b5:a2)}));
  assign y14 = {4{{1{p14}}}};
  assign y15 = (((!p2)&(^p5))|((p5<=p6)&(~p3)));
  assign y16 = (b3?b2:b0);
  assign y17 = ((b4?b0:b0)|(b3?a0:p15));
endmodule
