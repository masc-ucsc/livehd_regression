module expression_00737(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({{(-2'sd1),(-5'sd3)}}-{(5'sd6),(-3'sd1),(2'd3)})-(2'd3));
  localparam [4:0] p1 = {1{((3'sd0)>>>{2{((3'd5)^~(-4'sd2))}})}};
  localparam [5:0] p2 = {3{(2'd0)}};
  localparam signed [3:0] p3 = (((5'd29)==(5'sd11))!=={(5'd6)});
  localparam signed [4:0] p4 = (~&(2'sd0));
  localparam signed [5:0] p5 = (!(-3'sd0));
  localparam [3:0] p6 = {4{(-5'sd14)}};
  localparam [4:0] p7 = (~|{(~{(!(|{3{(3'd6)}})),(((4'd12)?(4'sd4):(4'sd5))?(!(-5'sd6)):((5'd31)?(4'sd4):(-3'sd1)))})});
  localparam [5:0] p8 = (3'sd0);
  localparam signed [3:0] p9 = (4'd0);
  localparam signed [4:0] p10 = (((3'sd2)?(2'sd1):(2'd2))|(~&{((-2'sd0)==(2'sd0))}));
  localparam signed [5:0] p11 = ((4'd1)==(-4'sd4));
  localparam [3:0] p12 = ({4{(2'd2)}}||(~|{2{(5'd6)}}));
  localparam [4:0] p13 = (+(((4'sd6)<=(-3'sd0))?((3'd1)?(5'sd15):(5'd15)):((3'sd0)?(-2'sd1):(5'd6))));
  localparam [5:0] p14 = {3{((-4'sd5)>=(2'sd0))}};
  localparam signed [3:0] p15 = (((4'sd2)?(-3'sd2):(4'd13))<(~&((4'sd7)?(5'd20):(3'd6))));
  localparam signed [4:0] p16 = {1{(((2'sd1)?(2'd3):(5'd23))?(~^(-(-2'sd1))):((4'd14)>>>(4'd8)))}};
  localparam signed [5:0] p17 = ((3'd0)?(-5'sd7):(3'sd3));

  assign y0 = (5'd21);
  assign y1 = (|{3{(a4?p11:b5)}});
  assign y2 = {1{((6'd2 * p6)&(p5==p16))}};
  assign y3 = {{{{{a2,a3,a5}},{b0,a0,b0}}},{{a4,a1},{p0,a2},{a3,b2}},{{{b5,a2,b3},{{p3,a0,b5}}}}};
  assign y4 = (((b5?b3:b3)<=(a0?b4:b2))-{{p2,p15,p16},{p12,p17,b3}});
  assign y5 = (|{(&(~{2{(~|(p5&p13))}})),{1{{3{(p10?p15:p7)}}}}});
  assign y6 = ((((~^b1)<<(p6+a4))>>((~a2)>>{p5,p3,b2}))<<<{{(&((~|(+p17))^~(a1^~p5)))}});
  assign y7 = {2{($unsigned({2{p12}}))}};
  assign y8 = (-a4);
  assign y9 = (&((a5>>>b3)-(b2<b3)));
  assign y10 = (((|(4'd8))!==(2'd1))===(&{3{(3'd4)}}));
  assign y11 = ((~p0)?$unsigned(p12):(a2+b1));
  assign y12 = (~&(p7>>>p8));
  assign y13 = (~((((-p12)&(3'sd2))<<<$signed(((b4))))&(4'd13)));
  assign y14 = (5'd18);
  assign y15 = (((b1&a0)<<(p13/a3))<<<(|((a1!==a4)!=(p0!=p14))));
  assign y16 = $unsigned(((a2&b5)&(p11?p6:a2)));
  assign y17 = {{{2{p16}},(a5&p10),(p14<<<a1)},{1{({4{p3}}==(b4<=p7))}},{{b2,p17,a3},(~^(~&b0))}};
endmodule
