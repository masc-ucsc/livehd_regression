module expression_00632(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(|(5'sd11))}?{(5'd12),(2'sd1),(2'd0)}:(~(2'd0)));
  localparam [4:0] p1 = {1{{4{{2{(2'sd0)}}}}}};
  localparam [5:0] p2 = {3{{2{(^(5'd12))}}}};
  localparam signed [3:0] p3 = ((&(~&(4'd6)))&((3'd0)?(4'sd0):(5'd21)));
  localparam signed [4:0] p4 = ((|(3'd7))<<<(+(-2'sd0)));
  localparam signed [5:0] p5 = (((3'd4)?(-2'sd0):(-4'sd7))?((2'sd0)?(-4'sd6):(-4'sd6)):((4'sd1)?(3'sd3):(4'd7)));
  localparam [3:0] p6 = (+((5'sd6)<<(-3'sd1)));
  localparam [4:0] p7 = (5'd25);
  localparam [5:0] p8 = ({(4'd7),(-2'sd0),(3'sd1)}<<<{(-4'sd2),(2'sd0),(3'd1)});
  localparam signed [3:0] p9 = ((((5'd21)>=(5'd6))!==((-3'sd3)?(4'd3):(3'sd3)))?((-2'sd0)?(3'sd3):(-3'sd3)):((2'd3)?(-3'sd0):(3'd0)));
  localparam signed [4:0] p10 = {4{(|(-(~^(5'd30))))}};
  localparam signed [5:0] p11 = (-5'sd2);
  localparam [3:0] p12 = (((5'd8)?(5'sd10):(4'd5))-((-3'sd1)<(-2'sd0)));
  localparam [4:0] p13 = ((&{(((3'sd3)<<(-3'sd3))>>{(4'sd4),(4'd13)})})==(((-3'sd0)>>>(5'sd8))?((-3'sd0)!=(-2'sd0)):(-{(-4'sd2)})));
  localparam [5:0] p14 = {{4{(4'd2)}},{{(3'd4),(-2'sd1),(5'd22)}},{1{{3{(3'd5)}}}}};
  localparam signed [3:0] p15 = (-3'sd2);
  localparam signed [4:0] p16 = ((((5'd12)-(5'd5))==(^((-3'sd0)!==(-5'sd15))))!==(((2'd1)>=(4'd12))||(4'd2 * (5'd11))));
  localparam signed [5:0] p17 = (~^((4'd2 * (-(4'd8)))>{(5'd8),(4'd5),(5'sd13)}));

  assign y0 = {1{{3{(+{3{a0}})}}}};
  assign y1 = ({(~&p6),(~&p0)}|((p9-p2)>>>{4{p6}}));
  assign y2 = (a4>p1);
  assign y3 = (~&({(5'd7)}==={(b3?b5:a2),(a0===b4)}));
  assign y4 = {4{(-{1{(~|a5)}})}};
  assign y5 = ((p15?p4:b3)<=$signed($unsigned(b4)));
  assign y6 = (^(p17^~p6));
  assign y7 = (+(+$signed(((a2?a5:b1)<<<(&{p0,b4,p7})))));
  assign y8 = ({({p11,p7,p13}<<$unsigned({p11,p10})),{((4'd2 * p1)>>$unsigned(p12)),{1{$unsigned({p13,p3,p3})}}}});
  assign y9 = ((3'd2)<<<{(a1!=p4),(a3<p15),{p17,b3,p10}});
  assign y10 = ({3{(p14&&p16)}}^~(({2{a1}}===(a5+b0))-(&(p3&p11))));
  assign y11 = (-5'sd13);
  assign y12 = {4{(a5?p16:b3)}};
  assign y13 = (b4?p15:b1);
  assign y14 = (5'd2 * (a2&&a1));
  assign y15 = (~&{4{(^b0)}});
  assign y16 = (&p13);
  assign y17 = (2'sd1);
endmodule
