module expression_00893(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(3'sd3),(5'd21)};
  localparam [4:0] p1 = ((({1{(2'sd1)}}==={2{(2'd3)}})|({4{(5'd27)}}||((3'sd3)|(-2'sd1))))===({1{((3'd4)<<<(-5'sd3))}}<=(((-2'sd0)||(3'sd2))&((3'sd1)>(4'd11)))));
  localparam [5:0] p2 = ((5'sd8)>=(-(((-4'sd6)>>(3'd6))==(&(-3'sd0)))));
  localparam signed [3:0] p3 = (+(+{3{(!(&(3'd6)))}}));
  localparam signed [4:0] p4 = (6'd2 * (5'd15));
  localparam signed [5:0] p5 = ((((4'sd7)?(4'd8):(4'd7))/(5'd11))?(&(((2'sd1)<=(-4'sd0))!=(~(4'd6)))):(~^(((3'sd3)?(2'd1):(-4'sd3))==(4'd2 * (3'd2)))));
  localparam [3:0] p6 = {(6'd2 * (+(2'd2))),(+((3'd6)-(3'd1))),({(4'sd6)}>{(-4'sd5)})};
  localparam [4:0] p7 = (&((~^(~^(-2'sd0)))?((3'd1)?(5'd21):(5'd1)):(|((4'd0)?(4'd10):(5'sd15)))));
  localparam [5:0] p8 = ((-5'sd1)-(-{3{((-4'sd3)<<<(2'd0))}}));
  localparam signed [3:0] p9 = ((&{(3'd0),(-4'sd5),(2'sd0)})+({(3'sd3),(4'sd7),(5'd16)}>>>((2'd2)>=(5'd2))));
  localparam signed [4:0] p10 = ((3'd3)==(-5'sd6));
  localparam signed [5:0] p11 = ({(-2'sd1)}^((5'd22)<<<(2'd2)));
  localparam [3:0] p12 = ((((5'd19)>(4'd3))^(^((-5'sd8)<(-2'sd1))))!==(&(|(((2'sd1)?(4'd15):(-3'sd0))<<{(4'd14),(-3'sd1)}))));
  localparam [4:0] p13 = ((((2'sd0)?(2'sd0):(3'd5))^~((4'd15)>>(5'd26)))+((-2'sd1)?(-3'sd3):(5'd17)));
  localparam [5:0] p14 = ((5'd22)?(3'd1):(3'sd2));
  localparam signed [3:0] p15 = {3{(-(^(5'd28)))}};
  localparam signed [4:0] p16 = ((3'd3)?(4'd7):(-3'sd1));
  localparam signed [5:0] p17 = {4{((5'd12)===(-5'sd13))}};

  assign y0 = (~((|(~&(3'd0)))&(^(-2'sd0))));
  assign y1 = {2{{p10,p13,p15}}};
  assign y2 = (((p15<<p1)?(p16<=p6):(a1!==b1))!={(p8?p3:b2),(p16&a2)});
  assign y3 = (b1<<b1);
  assign y4 = (^(+((~(+{4{(+p10)}}))||(((b3===a4))?(a1?p16:p8):{1{(a5>a5)}}))));
  assign y5 = ((p9?p16:p4)?(a4!==a2):(p13?p6:a5));
  assign y6 = (~^(~((&(p12<p8))/b0)));
  assign y7 = (~^((!(b1?b1:a2))===((5'd29)?(b4?a3:b5):(~&a3))));
  assign y8 = (3'd3);
  assign y9 = (~|(((p14&&p2)!=$signed((-a0)))&&((p1<<a1)>{a0,a3,b4})));
  assign y10 = {{((a0===b0)!==(a1<<b2))}};
  assign y11 = {(~(|a2)),{b1,p17,p4}};
  assign y12 = {2{(-4'sd6)}};
  assign y13 = ((a2?a5:b0)||(b1*a3));
  assign y14 = (((4'd9)>>((p12*p4)+(3'd4)))>>>((+$unsigned((p10>>p0)))<<(+((p7!=p1)))));
  assign y15 = (&(-(((a4===b5)!==(~^b3))?((&b0)>=(4'd2 * a2)):((a2&&b1)||(b1!=a2)))));
  assign y16 = (b1==p8);
  assign y17 = ((b1?p1:b2)?(p16?p13:p6):(p11?b5:p4));
endmodule
