module expression_00739(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(&((~|((2'd1)?(4'd13):(4'd9)))?{(~|(~(3'd0)))}:((3'd1)?(3'd0):(2'd3))))};
  localparam [4:0] p1 = (((((4'd12)^(4'sd4))==(6'd2 * (5'd23)))&&(((5'sd5)/(5'd27))>=((2'sd0)^~(3'd6))))<<(5'd2 * ((2'd3)-(3'd5))));
  localparam [5:0] p2 = (~^(~((5'd22)<<<(4'sd1))));
  localparam signed [3:0] p3 = {(((5'sd13)&(-4'sd3))>{(-4'sd3),(-4'sd0),(3'sd0)}),(((4'sd6)>=(2'd1))!==((4'd7)?(2'd1):(2'd1))),((^(3'd6))!=((5'd3)==(5'd22)))};
  localparam signed [4:0] p4 = (!({(4'sd6),(2'd1)}-(~&(5'sd9))));
  localparam signed [5:0] p5 = {{(5'sd12),(2'd0),(5'd17)},((3'sd2)^(4'sd6)),{(5'd28),(2'd3),(5'd12)}};
  localparam [3:0] p6 = ({4{(3'd0)}}<<<(^(4'd7)));
  localparam [4:0] p7 = (-3'sd1);
  localparam [5:0] p8 = (6'd2 * ((4'd9)>=(5'd16)));
  localparam signed [3:0] p9 = (5'd22);
  localparam signed [4:0] p10 = {(5'sd1)};
  localparam signed [5:0] p11 = (~&{1{((&{2{((-2'sd1)^~(2'd1))}})>{3{((2'd3)>>(2'd2))}})}});
  localparam [3:0] p12 = {4{((!(4'sd5))<<(^(2'd0)))}};
  localparam [4:0] p13 = ((((4'sd7)?(2'sd1):(-5'sd0))?{(5'd5),(4'sd6)}:{1{(2'd1)}})?{((2'sd1)?(-2'sd1):(3'd2)),((5'sd14)?(4'd1):(-5'sd4))}:{3{(!(4'sd5))}});
  localparam [5:0] p14 = ((-(+(-(2'sd0))))===(4'd1));
  localparam signed [3:0] p15 = (4'd3);
  localparam signed [4:0] p16 = (|(&((-4'sd6)|(-4'sd5))));
  localparam signed [5:0] p17 = (~^{4{(-2'sd1)}});

  assign y0 = (((b4?b1:b4)==={{1{{a4,a3,a5}}}})||((b5?a5:a4)?{1{{3{b1}}}}:(a2?b3:a3)));
  assign y1 = (~^{1{{3{((~$unsigned((p10>=p6))))}}}});
  assign y2 = $signed(($signed({{{b2,a5}},$signed($unsigned({p5}))})>={(((-4'sd2)^~(b0!==b5))>=(2'd2))}));
  assign y3 = ($unsigned({3{b1}}));
  assign y4 = ({{3{p11}},{a0}}|((2'd1)-(p5<<p5)));
  assign y5 = ((2'd2)?(p6==p3):(p7>>>p2));
  assign y6 = (!{1{{2{(p14?p1:p15)}}}});
  assign y7 = (2'd2);
  assign y8 = (&(!{($unsigned(((p9)!=(&a5)))^~(-{(~|a5),{a0}}))}));
  assign y9 = ((a4?b5:a5)*(b5|a0));
  assign y10 = (2'd3);
  assign y11 = (~(&((((a4/p6)/p14))!=(2'sd0))));
  assign y12 = {3{({2{p0}}<<{2{p8}})}};
  assign y13 = (((b0===b3)&{a5,b2,b5})>=$unsigned(((3'd2))));
  assign y14 = (4'd1);
  assign y15 = ((4'd2 * a1)^~{b4,b1});
  assign y16 = {((~^(+((p11)>>(a2))))|$signed(({2{p8}}<<<((&b2)))))};
  assign y17 = (p5^p12);
endmodule
