module expression_00069(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{3{(4'sd7)}},((2'd3)>>(2'd0)),{(-2'sd1),(5'sd14)}};
  localparam [4:0] p1 = {3{(&(2'd0))}};
  localparam [5:0] p2 = ({{{(-3'sd1)},{1{(5'd3)}},{4{(-4'sd5)}}}}>=(((-4'sd5)^(4'd0))<=((4'd11)===(2'sd1))));
  localparam signed [3:0] p3 = (^(((-3'sd0)>(-3'sd2))<={(3'sd2),(5'd20),(-5'sd14)}));
  localparam signed [4:0] p4 = ({4{(2'd3)}}<<<{1{(2'd3)}});
  localparam signed [5:0] p5 = ((5'sd2)?(-5'sd4):(3'd7));
  localparam [3:0] p6 = (5'd11);
  localparam [4:0] p7 = ((4'd4)>>(-5'sd1));
  localparam [5:0] p8 = (2'd1);
  localparam signed [3:0] p9 = ((((-2'sd1)>=(-4'sd7))<=((3'd6)==(3'd3)))===(~|(((5'd7)<=(5'd3))?((5'd19)>(2'd1)):((-5'sd15)?(2'd3):(-2'sd0)))));
  localparam signed [4:0] p10 = ((3'd2)&(5'd9));
  localparam signed [5:0] p11 = (3'd5);
  localparam [3:0] p12 = {((2'd0)?(2'd1):(5'd19)),((-5'sd9)?(3'd6):(-2'sd1))};
  localparam [4:0] p13 = (((~|(3'd4))||(+(5'sd8)))<=(&(~(-(!(-5'sd2))))));
  localparam [5:0] p14 = ({(-4'sd3)}?{(5'd0)}:{(-3'sd0),(4'd3),(-5'sd13)});
  localparam signed [3:0] p15 = {3{({4{(2'sd0)}}?(-(-2'sd1)):((-4'sd0)<(2'sd1)))}};
  localparam signed [4:0] p16 = {1{(|{3{{3{(5'sd9)}}}})}};
  localparam signed [5:0] p17 = {(|(!(((-3'sd1)?(2'sd1):(-3'sd2))?((3'd2)||(5'd1)):((3'sd0)<<(2'sd1)))))};

  assign y0 = {4{(a0==b2)}};
  assign y1 = (6'd2 * (2'd3));
  assign y2 = (((a0?p17:a3)?(p6?b4:b5):(!p8))&&((~&(|a5))>(~&{4{a5}})));
  assign y3 = {1{((^(-3'sd0))?((p11?a0:a0)):{2{(2'd2)}})}};
  assign y4 = {{p1},(p4?a3:p16),{a4}};
  assign y5 = ($unsigned((((p2*p10)^(p14-p4))^((p0&p13)==$unsigned(p16))))+(((p4%p0)==(p0==p5))<((p7-p3)>(p14*p2))));
  assign y6 = (((!(p10-p7))==(~|(p15^p1)))|((^{4{p2}})&&(~|(p15&p1))));
  assign y7 = (4'sd4);
  assign y8 = (3'd7);
  assign y9 = (!(!(-2'sd1)));
  assign y10 = ((p17?b4:p9)+$unsigned(({4{a3}})));
  assign y11 = (b1|p14);
  assign y12 = (~|(~|(4'd15)));
  assign y13 = (a2>b1);
  assign y14 = ((($unsigned($unsigned(p10))&&(p14||p15)))>((a0&&b4)===(b2^~a5)));
  assign y15 = ({(5'sd11),(p12<<<p17)}&((2'sd1)|(5'd26)));
  assign y16 = {((b1+b2)?(a4?a1:p17):(5'sd14)),{{a4,a4},(4'sd2)}};
  assign y17 = {((+(!(~{$signed((|{p7,p4,a3}))})))<<<((a5?a2:b1)?{p6,b5,b4}:(a3!==b3)))};
endmodule
