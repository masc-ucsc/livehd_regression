module expression_00987(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((!(4'sd2))*(4'd15));
  localparam [4:0] p1 = {(((3'd3)<(-5'sd9))+{(5'sd11),(3'd7)}),{4{(3'd2)}},(&{(^(-2'sd0)),((-2'sd0)<=(-5'sd0))})};
  localparam [5:0] p2 = (~((3'sd2)>>>(~&(3'd7))));
  localparam signed [3:0] p3 = ({((3'sd2)!=(5'd16)),(!{(4'd3),(3'd4),(5'd12)})}^~((~((-5'sd12)+(5'sd1)))>>(-{(2'd0),(5'sd0),(-2'sd1)})));
  localparam signed [4:0] p4 = {3{(4'd5)}};
  localparam signed [5:0] p5 = (+{2{(4'sd4)}});
  localparam [3:0] p6 = {3{{(3'sd0),(3'sd1),(5'sd12)}}};
  localparam [4:0] p7 = (~^(((+(3'd3))<=((3'sd2)?(5'd9):(-2'sd0)))!={(((4'd13)?(3'd7):(-3'sd0))&((-2'sd1)?(-5'sd10):(3'sd0)))}));
  localparam [5:0] p8 = {{((2'sd1)?(3'sd3):(3'sd0)),{(3'd7)},(&(3'sd2))},{{(5'd22),(3'sd0),(-3'sd2)},((-3'sd3)>(-2'sd1)),{(4'sd3)}}};
  localparam signed [3:0] p9 = {({(~|(3'd7)),((4'd14)?(-3'sd0):(2'sd1))}?((5'sd4)?(-3'sd2):(5'sd4)):(!(~&((4'd9)?(3'd2):(3'd1)))))};
  localparam signed [4:0] p10 = (|(-2'sd1));
  localparam signed [5:0] p11 = {((~&(-2'sd1))?{(5'sd7)}:(-4'sd4)),(+({(2'd3),(3'sd2),(5'd14)}===(2'd3))),(&(^((2'd2)?(2'd1):(5'd25))))};
  localparam [3:0] p12 = ((((-5'sd5)>=(4'd5))>=((-5'sd9)?(-2'sd1):(2'sd1)))>((~|(5'd14))|((-3'sd0)?(-4'sd4):(3'd4))));
  localparam [4:0] p13 = (~&((-2'sd1)?(2'sd1):(4'd1)));
  localparam [5:0] p14 = (((-2'sd1)&&(5'd29))?{(-2'sd0),(3'sd2),(2'd2)}:{(2'd1),(2'sd0)});
  localparam signed [3:0] p15 = (((3'sd1)||(-4'sd1))<<((-4'sd4)>(2'sd0)));
  localparam signed [4:0] p16 = ((((5'sd1)===(3'd0))+(2'sd0))^~{4{(4'd13)}});
  localparam signed [5:0] p17 = (~{3{(-5'sd12)}});

  assign y0 = ($unsigned($unsigned(((b4?a2:b5)==(-p11))))!=((-5'sd9)?(p10):{b3,b5,b4}));
  assign y1 = (((~(a2==b2))&(|(-p17)))|((5'd2 * a0)?(p1|a2):(a3%b3)));
  assign y2 = ((-2'sd1)!=={2{(a4+b5)}});
  assign y3 = (((p12-p4)?{2{p2}}:(b5?a0:p11))>={3{{p6}}});
  assign y4 = ((((p17<<p5)>=(p8>>>p13))>>(4'd2 * (p13||p1)))>=(5'd2 * {a2,b0,p8}));
  assign y5 = {p2,p6};
  assign y6 = (~^(&{(~|(~^b1)),(|(~^a1)),{a3,b3}}));
  assign y7 = {{1{(|(+{p7,a3,a4}))}}};
  assign y8 = {((-5'sd2)&$unsigned((a1^p11)))};
  assign y9 = {3{p12}};
  assign y10 = ((p9?p6:p14)?(~p13):(p8?a2:p8));
  assign y11 = (({1{(^p16)}}!=(a2!==b5))>=((a0||a1)?(^b4):(+a1)));
  assign y12 = {(a0|a2)};
  assign y13 = ((b2?b5:a3)?(b1?a1:a0):(b0?a3:p12));
  assign y14 = (~^({(~|p11),(p14?p4:p5)}?(p6?p6:p6):(|(a2?p16:p11))));
  assign y15 = (((p8*a5)==(a2?b3:a5))<((a4?b5:a5)&(b5+a4)));
  assign y16 = {{2{(a5>>b1)}},((a3||p3)-{b1,a5,a1})};
  assign y17 = $signed((~|((5'sd5)&((~b2)!==(a2<=b2)))));
endmodule
