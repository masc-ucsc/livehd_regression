module expression_00046(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'd2 * (~^((4'd7)>=(5'd16))));
  localparam [4:0] p1 = {1{{1{{4{{3{(3'd2)}}}}}}}};
  localparam [5:0] p2 = ((2'sd1)?((4'd1)?(3'sd2):(3'd0)):(5'd1));
  localparam signed [3:0] p3 = {1{({1{{4{(5'sd10)}}}}^~{3{(3'sd3)}})}};
  localparam signed [4:0] p4 = (^(~&(|((((-5'sd8)?(3'd7):(-5'sd4))&((5'sd6)%(5'd11)))<<(((3'd5)*(3'd0))<((5'd6)?(-4'sd1):(5'sd0)))))));
  localparam signed [5:0] p5 = (({2{(5'sd1)}}?(-(-2'sd1)):((4'd3)?(5'd15):(3'd7)))!=(((3'd4)&(4'd1))?((-4'sd0)?(4'd5):(2'sd0)):{1{(4'sd4)}}));
  localparam [3:0] p6 = ({3{(2'd3)}}?(|(|{3{(2'sd0)}})):(-((2'd3)?(3'd7):(4'd9))));
  localparam [4:0] p7 = (((6'd2 * (2'd2))+{2{(-5'sd8)}})<<<(((4'sd5)?(2'd0):(3'sd2))&((3'sd1)<(2'd3))));
  localparam [5:0] p8 = ((~^((3'sd3)!==(5'd8)))!=((5'd28)?(4'd13):(4'd7)));
  localparam signed [3:0] p9 = ((&((3'd0)!==(-3'sd2)))!=={((4'd2)!=(2'sd0))});
  localparam signed [4:0] p10 = ((3'd0)%(3'd4));
  localparam signed [5:0] p11 = ((((5'd13)==(2'd2))?((5'd22)?(3'd5):(4'd10)):((3'd3)?(3'd2):(3'd2)))-(((4'd2)>>(2'd3))?((-4'sd3)%(3'd0)):((-2'sd0)+(4'd14))));
  localparam [3:0] p12 = ({(-4'sd5),(-5'sd5),(3'd5)}!=((3'sd1)?(2'd1):(2'd3)));
  localparam [4:0] p13 = ((-2'sd0)?(2'sd1):(2'sd0));
  localparam [5:0] p14 = (-(4'd10));
  localparam signed [3:0] p15 = {2{{2{{2{(2'd3)}}}}}};
  localparam signed [4:0] p16 = ({(-3'sd3),(-2'sd1),(-5'sd4)}=={(5'sd0),(3'sd1)});
  localparam signed [5:0] p17 = ({2{(&(4'sd3))}}<<({3{(-2'sd1)}}^((5'sd15)?(5'd7):(-4'sd0))));

  assign y0 = (!(3'd5));
  assign y1 = (({1{p4}}=={p13,p16,p15})<<$signed({2{p5}}));
  assign y2 = (-2'sd0);
  assign y3 = ({3{p17}}?$unsigned((~^$signed(p8))):$unsigned((~^(b5===a0))));
  assign y4 = ({1{((p17?p4:a1)?(p13^p2):(p1?p11:b4))}}>>>(((p1-p9))?{p14,p1}:(p13!=p1)));
  assign y5 = (~&($signed($unsigned(a2))|(-2'sd0)));
  assign y6 = {2{{b1,p14,b0}}};
  assign y7 = ((~^(|(&{3{a4}})))?({3{p8}}?(-2'sd1):(~^b0)):(~|{3{(&a0)}}));
  assign y8 = (((a4<p12)!=(p1%p8))^~(-3'sd0));
  assign y9 = (5'd19);
  assign y10 = (p3>=p14);
  assign y11 = (-2'sd0);
  assign y12 = {4{a0}};
  assign y13 = (a2<<b0);
  assign y14 = {2{({1{(p3<=p6)}}?(+{2{p6}}):(p2?b2:p12))}};
  assign y15 = {$unsigned((4'sd1)),(a5<b1),$signed((~b1))};
  assign y16 = ((($signed(a3)?(2'd0):$signed(b3)))?((5'sd6)?(a2<a3):(a1?a3:p6)):(((-3'sd2)?(b4%a0):(b3?b1:b2))));
  assign y17 = (^{((a0>=p7)<<<(p7<<<p1))});
endmodule
