module expression_00798(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(~(!(-4'sd1)))}};
  localparam [4:0] p1 = (~^{1{(~^((-({2{(5'd12)}}>>((2'd2)>(4'd15))))!==(((-4'sd1)-(5'd25))?((4'd14)&&(3'd5)):((5'd18)+(5'd14)))))}});
  localparam [5:0] p2 = ((2'sd1)-(4'sd2));
  localparam signed [3:0] p3 = (+((3'd6)>>(5'd26)));
  localparam signed [4:0] p4 = (|((+(5'sd4))||((3'd4)<<<(5'd26))));
  localparam signed [5:0] p5 = ((5'sd9)<<<(3'd6));
  localparam [3:0] p6 = {(~&{(3'd6),(2'd2),(2'd0)}),(~|{(-4'sd3),(3'sd2)}),(~&(&(3'd1)))};
  localparam [4:0] p7 = ((((6'd2 * (2'd0))!==(4'd2 * (3'd5)))>>>((4'd2 * (5'd25))+((5'd26)>(5'd4))))-((((3'sd3)||(2'sd1))&((3'd0)/(5'd9)))<(((3'sd0)!=(-2'sd1))|((-4'sd1)|(4'sd6)))));
  localparam [5:0] p8 = ((2'd3)<=(5'd16));
  localparam signed [3:0] p9 = ({1{(-3'sd1)}}!==(3'd4));
  localparam signed [4:0] p10 = ((((2'd2)||(-5'sd12))!==((3'd0)*(4'd4)))==(((2'd3)/(-4'sd6))<<<((-4'sd5)==(2'sd0))));
  localparam signed [5:0] p11 = (4'd11);
  localparam [3:0] p12 = (5'd13);
  localparam [4:0] p13 = (-((|((3'd2)===(2'sd1)))==(2'd3)));
  localparam [5:0] p14 = ({(5'd8),(-3'sd2),(-5'sd9)}<<(!{1{{(-3'sd2),(2'd2)}}}));
  localparam signed [3:0] p15 = ((|{3{(~|(4'd7))}})>(&(|{2{(~^(2'd2))}})));
  localparam signed [4:0] p16 = (+(3'sd3));
  localparam signed [5:0] p17 = ((!(~{3{(3'sd0)}}))?(!(&(^(4'd13)))):((2'd3)?(2'd2):(2'sd0)));

  assign y0 = {{4{(-p16)}},{{b1,p15},(p4?a5:a0)},((~^p11)?(^p14):(p12?p7:a4))};
  assign y1 = (5'd13);
  assign y2 = ((b0?p10:p3)?(p1?p13:p6):(3'd2));
  assign y3 = (4'sd1);
  assign y4 = (-3'sd2);
  assign y5 = (3'd1);
  assign y6 = (5'sd0);
  assign y7 = ((((b2?p1:b0)<=(b2<p9))<=(p16?p6:p14))|(3'd2));
  assign y8 = (5'd20);
  assign y9 = ((~(b0*b3))/a5);
  assign y10 = (4'd9);
  assign y11 = (4'd2 * (a1|a2));
  assign y12 = (((|(p11?b0:a1))-{4{a1}})?((a0?b0:b3)>(a3^~b5)):({3{a1}}?(!b2):(b2!=b0)));
  assign y13 = {{(-4'sd6)},(&(^{p14,a0,b4}))};
  assign y14 = {3{{1{p6}}}};
  assign y15 = {2{{4{{2{p16}}}}}};
  assign y16 = {{{1{{3{p14}}}}},$signed((b5!==a4)),$signed({{2{b4}}})};
  assign y17 = {2{(4'd2)}};
endmodule
