module expression_00359(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!((-3'sd3)%(2'd0)));
  localparam [4:0] p1 = ({1{((-5'sd4)?(3'sd1):(-3'sd1))}}?{4{(5'd12)}}:(((-4'sd3)?(2'd3):(4'd10))?{1{(3'd7)}}:((2'd3)?(3'd3):(4'd12))));
  localparam [5:0] p2 = (2'sd0);
  localparam signed [3:0] p3 = (((2'd3)!=(-2'sd1))<=(!(5'sd13)));
  localparam signed [4:0] p4 = {(-(2'sd0))};
  localparam signed [5:0] p5 = ((~^{{(-3'sd3),(-5'sd8)},((-2'sd0)!=(5'd22)),{(-5'sd5),(2'd0)}})^{(!(|(~&(-(^(3'sd1))))))});
  localparam [3:0] p6 = {({(2'd0)}?((5'd16)?(4'd4):(3'sd3)):{4{(4'sd2)}}),{3{{(-3'sd3),(5'sd14)}}}};
  localparam [4:0] p7 = ((2'd3)?(5'd27):(2'sd0));
  localparam [5:0] p8 = ((2'd3)-(-4'sd6));
  localparam signed [3:0] p9 = (!(3'd5));
  localparam signed [4:0] p10 = (~^(4'sd7));
  localparam signed [5:0] p11 = {((~(^(-3'sd3)))===(~|{(4'd11),(5'd8)}))};
  localparam [3:0] p12 = (-((-(4'sd6))<=((5'sd8)>(-5'sd12))));
  localparam [4:0] p13 = (4'sd0);
  localparam [5:0] p14 = (3'd4);
  localparam signed [3:0] p15 = (+{({(4'sd3)}==={(4'd15),(-3'sd2),(-3'sd1)}),(((2'sd1)>>>(2'd1))-(~(3'sd2))),{(5'sd2),(-4'sd0),(5'd22)}});
  localparam signed [4:0] p16 = (((&(3'sd3))<=(|(4'd14)))>>(+(((5'sd9)===(2'd1))%(3'd6))));
  localparam signed [5:0] p17 = ((~(^(-2'sd1)))||{(5'd7),(2'sd0)});

  assign y0 = {2{(((b0>b4)===$signed(b0))<<($unsigned({3{p1}})))}};
  assign y1 = ((^(!(2'd2)))||{(-5'sd2),(+p12)});
  assign y2 = ((p4?p5:p0)|(p12+p7));
  assign y3 = {2{{2{a1}}}};
  assign y4 = {($signed((-3'sd1)))};
  assign y5 = (~^((2'sd0)^(|(p14>>p8))));
  assign y6 = $signed({2{(((^p15))>{4{b5}})}});
  assign y7 = {(~^{(+(p17>>a1))}),(~|((|p6)<<<{p10,p6,p13})),(|(^(^(~a3))))};
  assign y8 = {((~^((!(a0>a1))>>>{(b4&&b5)}))^(~{(((~$unsigned((&(a1<=a4))))))}))};
  assign y9 = ((&((|p12)<<<(|p4)))?((|p9)*(p10&a3)):(~&((p8<<p1)+(p3-p15))));
  assign y10 = {{b0,b4},{1{a5}}};
  assign y11 = (a2?p14:p12);
  assign y12 = ({(b4),(p0?b0:b0),(p14?p8:p5)}&(-{(b4?p17:p12),$unsigned((-3'sd1))}));
  assign y13 = (($unsigned(b2)>>(b4&&b5))<=((a4)^~$unsigned(b3)));
  assign y14 = (!(~^(((p10^b2)>=(p13|b0))^{(|p9),(+p7),(p17||p16)})));
  assign y15 = {3{(-(+{2{(|b2)}}))}};
  assign y16 = ((&(~&({(b1>>>b0)}===(&(!a2)))))|(5'd2 * $unsigned((~^p1))));
  assign y17 = (~^(~(~|({3{p5}}?({4{a0}}):(2'd3)))));
endmodule
