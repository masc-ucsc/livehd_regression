module expression_00240(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{((3'sd0)|(-4'sd1))}};
  localparam [4:0] p1 = ({4{(2'd3)}}?((^(3'd3))<=((3'd7)?(4'd14):(-2'sd0))):((~&(3'd4))=={3{(4'd11)}}));
  localparam [5:0] p2 = ((4'd3)?(5'd22):(3'd0));
  localparam signed [3:0] p3 = ((~^{(4'sd6),(2'd0),(-2'sd0)})<<<({(5'd14),(-2'sd1)}?{(5'd21),(-5'sd11),(4'sd6)}:(+(-3'sd0))));
  localparam signed [4:0] p4 = (!(2'd3));
  localparam signed [5:0] p5 = {3{((-4'sd6)<<<(-3'sd1))}};
  localparam [3:0] p6 = ((2'd2)+((4'd4)|(5'sd4)));
  localparam [4:0] p7 = ((5'd11)<<<(-2'sd1));
  localparam [5:0] p8 = (((-(4'd11))/(5'd3))>>>(2'sd0));
  localparam signed [3:0] p9 = ((|((-5'sd12)?(4'd1):(5'd29)))?((5'd16)?(4'sd4):(5'd24)):(+((2'd3)!==(-3'sd2))));
  localparam signed [4:0] p10 = {(!(~(^(2'd0)))),(((2'sd0)&&(3'sd2))|{(2'd2),(3'd3)}),(^(3'sd3))};
  localparam signed [5:0] p11 = {{3{{(4'sd1),(5'd15),(-5'sd3)}}}};
  localparam [3:0] p12 = ((4'd4)!==(-2'sd0));
  localparam [4:0] p13 = (-4'sd4);
  localparam [5:0] p14 = (5'd21);
  localparam signed [3:0] p15 = (4'sd2);
  localparam signed [4:0] p16 = ((&(2'sd0))?((-4'sd0)^(-2'sd1)):((-4'sd5)===(-3'sd1)));
  localparam signed [5:0] p17 = (4'd15);

  assign y0 = ({(p13?p11:b2),(p13-a0),(p13>p9)}^~((b2<a5)+(p6?p17:p3)));
  assign y1 = {{(b5!==a4)},$unsigned((a4||a0)),((b0!==b2)^{p13,b4,b1})};
  assign y2 = (^(2'd0));
  assign y3 = {(a1?a3:b4),((a3?b4:a0)<=(~&a1)),((+p4)&{b4,b0,p9})};
  assign y4 = (~(((-4'sd6)<=(p17>>>b3))!=(~((p10<=p10)&(p7<<<p3)))));
  assign y5 = ($signed((b5?b0:b4))?{4{a4}}:$unsigned((b3?b4:a0)));
  assign y6 = (((~&b0)?$unsigned(a3):(b5===b0))?{1{{1{(p7?p8:p1)}}}}:(|{2{(~b0)}}));
  assign y7 = (((b1>=p15)*(a1<<<p7))?((p1?p12:a5)>>>(a5-a5)):((p11<=a1)<<<(b0!==a0)));
  assign y8 = (~|$unsigned((|(|(~&$unsigned(((~|(~(p1?p7:p8)))?((p1?p0:p17)?(~^p2):(!p1)):(-$signed($signed($signed(p10)))))))))));
  assign y9 = {$signed((2'd0)),(2'sd1),(p14?b0:p5)};
  assign y10 = (((b3^a4)>>$signed(a2))?(~|(b3?a5:b3)):({a0,b4,a2}|(~^b0)));
  assign y11 = (3'd4);
  assign y12 = ((~$unsigned({2{(|b4)}}))&{2{(+(^b2))}});
  assign y13 = {{4{(p0>=p12)}},{4{(b2||b5)}},(&{1{{2{(b2&b2)}}}})};
  assign y14 = (({b0,b1,a0}||(5'sd0))!=(-3'sd3));
  assign y15 = (b3/a1);
  assign y16 = ($signed(b4)?{1{p5}}:$unsigned(b0));
  assign y17 = ((6'd2 * (p0||p0))<({(p4<<p10)}^~(p12-p15)));
endmodule
