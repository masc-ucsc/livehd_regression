module expression_00098(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^{(~({(5'd24),(3'd5),(-4'sd3)}<<<{4{(-2'sd1)}})),{3{{1{(2'd3)}}}}});
  localparam [4:0] p1 = ((4'd12)^~(-4'sd0));
  localparam [5:0] p2 = {((2'd1)<=(-3'sd2))};
  localparam signed [3:0] p3 = (5'd31);
  localparam signed [4:0] p4 = {(((-4'sd3)?(4'sd4):(4'sd5))>>>((2'd0)<<(4'd4))),(((5'd3)>(4'd11))^{2{(2'd1)}}),(((-5'sd8)|(2'sd0))-((4'd12)|(5'sd4)))};
  localparam signed [5:0] p5 = (((2'sd1)?(5'sd15):(3'sd0))?((5'sd9)?(-4'sd4):(-5'sd1)):((3'd2)?(-2'sd1):(3'd7)));
  localparam [3:0] p6 = (-3'sd3);
  localparam [4:0] p7 = {3{(-3'sd3)}};
  localparam [5:0] p8 = (2'd3);
  localparam signed [3:0] p9 = {4{(3'd6)}};
  localparam signed [4:0] p10 = ((((4'd4)<<<(4'sd7))-{1{(3'sd2)}})?({1{(5'd23)}}&(~&(2'd3))):(((2'sd0)<<<(2'sd0))&&((-3'sd0)+(5'd22))));
  localparam signed [5:0] p11 = ((((3'd0)!=(2'sd1))&&((5'd18)?(5'sd12):(5'sd11)))?(((2'sd1)>(2'sd0))===((2'd3)?(2'sd1):(-3'sd2))):({(4'd9)}>={(-5'sd8),(-4'sd7)}));
  localparam [3:0] p12 = ((5'd2 * ((5'd28)!=(3'd0)))>={1{(~|((2'sd1)-(4'sd3)))}});
  localparam [4:0] p13 = (~^(~|((+(((4'd13)&(3'd6))>>>(~(-4'sd6))))!=(~&(+(~&(-(5'sd8))))))));
  localparam [5:0] p14 = ((4'd2)?(4'sd7):(4'd10));
  localparam signed [3:0] p15 = {1{((3'd5)<(5'd28))}};
  localparam signed [4:0] p16 = {2{((5'sd7)?(-5'sd6):(2'd0))}};
  localparam signed [5:0] p17 = (|(!(((3'd1)?(-5'sd15):(-5'sd6))?((2'sd0)?(2'd3):(5'd27)):((4'd11)?(5'd10):(5'd7)))));

  assign y0 = (5'd2 * (b2|b0));
  assign y1 = (&($signed(((~^p11)<<(!p5)))<=((~p0)||(p12||p5))));
  assign y2 = {(b4?a3:b0),(a0?p8:a3),(4'd1)};
  assign y3 = ((p17&&p5)?{p14,p12}:(p13<<<p2));
  assign y4 = (5'd14);
  assign y5 = (((p13!=b5)?$signed(p11):{p0,p12})+((p7>>>b0)>(p17^p7)));
  assign y6 = (~&{(&((+p14)^{p5,p7})),(!((^p15)+(p17==p14)))});
  assign y7 = {4{(^{2{a1}})}};
  assign y8 = (2'sd0);
  assign y9 = ((3'd6)*(p8?b1:b2));
  assign y10 = ({(a2?a1:b5),(|(a0|b0)),(a1?b4:b4)}===((b2?a2:b0)?{b4,b1,a0}:(b1||a5)));
  assign y11 = (~&{((p5<<<b5)|(b2&&a4))});
  assign y12 = ((((a0>>>b1)^(!a5))-(~(a1?b1:a5)))===(((b2?a0:b0)*(a0|a2))>(~&(|(b0&&b1)))));
  assign y13 = (((b5<b0)<(+(b5>>a2)))<(!{1{{2{(b3!=a0)}}}}));
  assign y14 = (|{(~&$signed($signed((a4-a2)))),(-((4'd12)<(~&a2))),{{a1,b0},$unsigned(a4)}});
  assign y15 = ((+(~&(a0&&b1)))||$signed((p14<a1)));
  assign y16 = (5'sd7);
  assign y17 = (&(-4'sd2));
endmodule
