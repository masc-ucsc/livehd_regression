module expression_00175(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(^(-4'sd7)));
  localparam [4:0] p1 = ({4{(5'sd8)}}==((5'sd8)?(-2'sd1):(5'd23)));
  localparam [5:0] p2 = {3{((5'd27)!=(3'sd2))}};
  localparam signed [3:0] p3 = {1{(~&(~&{2{{((2'd3)?(-5'sd3):(5'd7)),{2{(-5'sd8)}}}}}))}};
  localparam signed [4:0] p4 = (~^(~|{((2'd3)>=(-5'sd14)),(~(3'd6)),{(5'd29)}}));
  localparam signed [5:0] p5 = (~(|(^(|(-(+(~(|(^(~&(+(-(~|(4'd4))))))))))))));
  localparam [3:0] p6 = ((((-2'sd1)?(-4'sd1):(-3'sd3))^~(~&(2'd2)))||((5'sd6)?(4'd5):(-4'sd2)));
  localparam [4:0] p7 = (2'sd1);
  localparam [5:0] p8 = (~&(4'd2 * (3'd3)));
  localparam signed [3:0] p9 = (~^(3'd6));
  localparam signed [4:0] p10 = {{(|((-4'sd4)==(3'd2))),{(5'd1),(3'sd0),(3'sd3)}},(((4'sd3)^(4'd8))>=(~^((5'sd2)|(-3'sd0))))};
  localparam signed [5:0] p11 = {3{(((3'sd1)>=(-4'sd3))&((3'd5)>>>(5'sd10)))}};
  localparam [3:0] p12 = ((5'sd14)?(4'sd3):(2'd2));
  localparam [4:0] p13 = {4{(~(5'd2))}};
  localparam [5:0] p14 = (-(|(-(((5'd0)>(2'd2))<=(~^((-2'sd1)>(4'd14)))))));
  localparam signed [3:0] p15 = ({1{(5'd21)}}?((3'd2)?(5'd27):(2'd1)):(^(3'd0)));
  localparam signed [4:0] p16 = (3'd5);
  localparam signed [5:0] p17 = (4'd12);

  assign y0 = {{(-5'sd15),(5'sd7),(5'd10)},(-2'sd1)};
  assign y1 = (~^((p2<p9)?{p8,p6,p8}:(p17>>p16)));
  assign y2 = (~^((((b2||p4)+(a1>>p0))<{3{a4}})>>(2'sd1)));
  assign y3 = {1{(~|{2{{1{{1{(|{2{{3{p9}}}})}}}}}})}};
  assign y4 = ($unsigned(p14)!=(a1));
  assign y5 = (&(({(p12+p9)}|(|{2{p9}}))<<<(~^((~|{p2,p2,p16})>>{4{p1}}))));
  assign y6 = {4{{3{b3}}}};
  assign y7 = {(~{(p2+a3)}),(~&{{a4,p1,p0}}),{p4,p15,p8}};
  assign y8 = (!{$signed({{p16},(-p17),{2{p3}}})});
  assign y9 = (&(-$unsigned(((~&p15)?$unsigned(b1):$unsigned(b2)))));
  assign y10 = $signed($unsigned((+$signed(((b1)!=={b1})))));
  assign y11 = ((~^(4'd14))>=(5'd3));
  assign y12 = (!((4'd4)&{2{b0}}));
  assign y13 = (~((+(~&((a3>>>a1)?(b5==p12):{b1,a4})))>=({(^b3),{p0,p1},(a2-b0)}&(5'sd4))));
  assign y14 = {1{(!(!p13))}};
  assign y15 = ((b3|a4)/p6);
  assign y16 = (~|(~|(|(((p8||p15)|(~^p13))?((a3==p12)||(p5!=p8)):(~|(a1?a0:p12))))));
  assign y17 = ((-({b3,b5}||(+a0)))!=={((a5?b1:a2)>(!a3))});
endmodule
