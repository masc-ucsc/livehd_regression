module expression_00821(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(4'd2 * (~|((5'd28)>(4'd6)))),(-((+((4'sd3)>=(2'sd0)))^(2'sd1)))};
  localparam [4:0] p1 = (^(+{((4'd15)?(-2'sd0):(5'd11))}));
  localparam [5:0] p2 = {((5'd25)+(2'd1)),((-2'sd1)?(5'd28):(3'd7)),((-3'sd0)>(3'd3))};
  localparam signed [3:0] p3 = {2{(~{(3'sd0),(-3'sd2)})}};
  localparam signed [4:0] p4 = (4'd9);
  localparam signed [5:0] p5 = (((!(4'd12))-((-5'sd11)<<(4'd7)))^(3'd5));
  localparam [3:0] p6 = ((-2'sd1)!==(4'd7));
  localparam [4:0] p7 = (~^({1{({2{(5'sd2)}}<=((2'd2)>=(5'd22)))}}!==(^((^((3'sd1)-(4'sd4)))<<((4'sd4)>>(2'd0))))));
  localparam [5:0] p8 = {(2'd3)};
  localparam signed [3:0] p9 = (~^(3'd1));
  localparam signed [4:0] p10 = ({((3'sd2)<<(5'd28)),(|(4'd4)),{(-2'sd0)}}>>>((2'd3)>>((5'd23)^(2'd1))));
  localparam signed [5:0] p11 = {(5'sd6),(-2'sd0),(-3'sd1)};
  localparam [3:0] p12 = {{{(-4'sd1),(-2'sd0)},{(3'sd3),(2'd0)},((-3'sd2)<<(4'sd0))},{{(2'd0),(-2'sd0),(2'd1)},{1{((-4'sd0)>(-5'sd8))}}}};
  localparam [4:0] p13 = (4'd1);
  localparam [5:0] p14 = (~|(-(&(((2'd3)?(-4'sd4):(-3'sd2))?{3{(5'sd14)}}:(((-4'sd0)&(-3'sd3))+(|(4'd0)))))));
  localparam signed [3:0] p15 = (3'd7);
  localparam signed [4:0] p16 = (2'd0);
  localparam signed [5:0] p17 = (|(5'd2 * (!(~^(4'd14)))));

  assign y0 = {4{b3}};
  assign y1 = (((a2^~b4)?(a4<<<p9):(p1>=a0))<=((5'd2 * a0)>>(p9?p1:b3)));
  assign y2 = (-((a2|p16)?(p4?p17:b2):$unsigned($signed(p16))));
  assign y3 = (({a5,b3,b4}>>>(b5^~b1))===({a4,b0,a5}||(a4&a0)));
  assign y4 = ((3'd5)<(4'sd3));
  assign y5 = (((p7^~p16)?(b0?b4:b5):(a5?p15:p12))<((!(b0?b2:a0))?(b3?p16:b0):(b1>>>b0)));
  assign y6 = {{4{a5}}};
  assign y7 = {{(a1>a2),{(a2||a2)},(a1^~p15)},(|(^((~^{p11,p9})|{a3,p2,p8})))};
  assign y8 = (&(4'sd6));
  assign y9 = {{3{{2{p14}}}},{{{(-5'sd6)}}}};
  assign y10 = $unsigned({$signed((|{(p4<<<a4),$unsigned(p7)})),{(~b0),(a4===a3),(b0)}});
  assign y11 = {((b5?a5:p6)?(p3-b3):(p15||b4))};
  assign y12 = (((&(a0|a0))===(+(|a4)))===((a4>b1)!=(~&(a0^a2))));
  assign y13 = (($signed((p12))<(p11>>>p11))|((p0-p5)^$unsigned($signed(p17))));
  assign y14 = (-4'sd2);
  assign y15 = (2'sd0);
  assign y16 = (((2'sd1)<((b4>>b5)!=(3'sd3)))<<{(a4?a4:b3),(3'sd1),(a0?b1:b2)});
  assign y17 = (~|$signed((~&{4{{2{p14}}}})));
endmodule
