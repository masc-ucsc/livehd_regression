module expression_00520(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'sd1)+(2'd0))-(3'd2))>>>{4{{2{(2'd1)}}}});
  localparam [4:0] p1 = {4{((5'd10)^(5'd3))}};
  localparam [5:0] p2 = (+(~(~^(2'sd0))));
  localparam signed [3:0] p3 = (-3'sd2);
  localparam signed [4:0] p4 = ({1{((4'sd1)!==(2'd1))}}|((3'd5)>>(-3'sd1)));
  localparam signed [5:0] p5 = (&(^(3'd0)));
  localparam [3:0] p6 = (~(&{(5'd27),(((3'd7)<(-5'sd14))<<<{(-2'sd1),(-2'sd0)})}));
  localparam [4:0] p7 = {(((-3'sd2)?(-2'sd1):(2'd3))<((5'd1)?(5'd21):(3'd1)))};
  localparam [5:0] p8 = {(5'sd1),(3'd4),(4'd1)};
  localparam signed [3:0] p9 = ({{2{(3'd4)}}}^~({(5'sd14),(4'd7),(3'd4)}-(((-4'sd2)>>(4'd2))+(|(-3'sd3)))));
  localparam signed [4:0] p10 = (~|{(+(((4'd2)<<(4'sd7))<<<(-(4'd10)))),(!({(-3'sd0)}!=(~(4'sd3)))),(~&((|(-2'sd1))<<<(4'd2 * (5'd19))))});
  localparam signed [5:0] p11 = (~^(^{({3{{2{(2'd0)}}}}>>{(+(2'd1)),{(2'd3)},(+(4'd12))})}));
  localparam [3:0] p12 = (~&({((2'd3)<=(3'd3))}&&{(4'sd7),(2'd1),(4'd12)}));
  localparam [4:0] p13 = (|(-2'sd0));
  localparam [5:0] p14 = (((2'd3)?(5'd26):(4'd1))?({1{(2'd0)}}|(+(2'd2))):(-2'sd1));
  localparam signed [3:0] p15 = (&((!((2'd3)>(4'd1)))*(!(^(-3'sd3)))));
  localparam signed [4:0] p16 = ((-5'sd12)^~(-5'sd7));
  localparam signed [5:0] p17 = {4{{2{(4'd2 * (2'd1))}}}};

  assign y0 = (((a5>>b3)<<<(~|(b0>=b3)))!==(+(~|($unsigned(b5)>>>(~^a1)))));
  assign y1 = {2{$signed(({b3,a3,a1}?$signed($unsigned(b1)):$signed($signed(a3))))}};
  assign y2 = (~(~^((p1?a3:p6)?{3{p8}}:(p14<p1))));
  assign y3 = (!{(|{(a3<<p6),(a2^a2)})});
  assign y4 = (~p14);
  assign y5 = (-2'sd0);
  assign y6 = (!{4{(&{3{p5}})}});
  assign y7 = {(5'sd3)};
  assign y8 = {((~^$unsigned(((2'sd1)>=(4'd12))))+(((~&a0)<=(~^p6))+(4'd2)))};
  assign y9 = $signed({{2{(({b4,a3})==={{b3,a0,a0}})}}});
  assign y10 = (~|$unsigned((!$unsigned((({b5,p16}&&(p5-a4))==({(-b4),{p4,a4,b3}}))))));
  assign y11 = (|{b2,b2});
  assign y12 = {{(a2===b4),(a1||p17),{b5}},$unsigned((&({3{a4}}==={b2,b4})))};
  assign y13 = (((~^(4'd7))>>$signed((p7>>p6)))^~((2'd1)&&((p17>=p1)>=(-p10))));
  assign y14 = ($signed(({(b3>>>a0),(b3&p2),(a0^~a4)}))-({(b1<=p11),{p9}}^~((p3^~b0)==(4'd2 * b0))));
  assign y15 = (3'd3);
  assign y16 = {2{(-2'sd1)}};
  assign y17 = (~(+((3'sd2)!=((4'd11)<<<(4'd11)))));
endmodule
