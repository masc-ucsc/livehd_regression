module expression_00334(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-4'sd7)===(-2'sd0))?((-3'sd2)|(4'd3)):{(3'd7)});
  localparam [4:0] p1 = (({(3'd2),(-5'sd2),(5'd19)}>>>(~|(5'd23)))+(~(~((5'd4)^(-2'sd0)))));
  localparam [5:0] p2 = (^(((5'd8)?(-5'sd15):(4'sd6))?(~^((5'd28)?(2'd2):(4'd7))):(4'd2 * (2'd2))));
  localparam signed [3:0] p3 = {({(|(-5'sd12)),{(2'd2)},{4{(-3'sd1)}}}-({(-5'sd12),(-4'sd6),(-3'sd2)}?(|(2'd0)):{(5'd20),(3'sd3),(2'd1)}))};
  localparam signed [4:0] p4 = ((~(&(((2'd1)&&(-3'sd3))!==((4'd5)<<(-3'sd1)))))-(((4'd0)!=(2'd3))||((3'd5)!==(3'd6))));
  localparam signed [5:0] p5 = (~{1{{(|({4{(4'd15)}}?{(2'd1),(-2'sd1)}:{3{(3'sd2)}})),(&(^(+((5'd11)?(5'sd4):(-2'sd1)))))}}});
  localparam [3:0] p6 = ((((3'd2)^~(4'sd3))&((5'sd13)>=(2'd2)))>>(((2'sd0)>(5'd9))>>>((3'sd3)&&(2'd0))));
  localparam [4:0] p7 = ((5'sd10)>>(5'd26));
  localparam [5:0] p8 = (3'd5);
  localparam signed [3:0] p9 = (~{3{{2{(3'd3)}}}});
  localparam signed [4:0] p10 = ((^{(4'd13),(5'sd11),(-2'sd0)})&((3'sd2)==(2'sd1)));
  localparam signed [5:0] p11 = ((~^(2'd1))?((2'sd1)?(-4'sd1):(5'sd4)):(3'd1));
  localparam [3:0] p12 = (4'd3);
  localparam [4:0] p13 = (|(3'd0));
  localparam [5:0] p14 = (|{4{(!{3{(2'd2)}})}});
  localparam signed [3:0] p15 = (5'd28);
  localparam signed [4:0] p16 = (-4'sd6);
  localparam signed [5:0] p17 = ((5'sd4)&&(-5'sd5));

  assign y0 = ({4{(p1?b0:p0)}}?{1{{3{(~&a5)}}}}:({3{p5}}?(b0?p10:p13):(~|b1)));
  assign y1 = (({(4'd2 * p13),(b3!==a0)}&&((b5^~p8)-$unsigned($signed(b2)))));
  assign y2 = (((~&b3)===(a4>=a1))&&{b4,p15,p8});
  assign y3 = (((p1/p13)?(3'd3):(p15>>>p11))?((p8?p10:p17)?(p8||p4):(p16?p9:p3)):((p7^p5)!=(4'sd5)));
  assign y4 = (^(((+(|a5))<<((^p17)))<=((a3===a0)>(+(b2===a5)))));
  assign y5 = {3{p14}};
  assign y6 = (&((~^({p10,b4}?(b1+p1):(|p17)))?((!p8)?{p10,p9,p9}:(~&a2)):(~((~^p3)!=(b1===b4)))));
  assign y7 = ((!$signed((-2'sd0))));
  assign y8 = ((a1?a5:b3)||(p11>>b0));
  assign y9 = ({3{{1{p16}}}}<<<({1{(~p14)}}==(p0<<p6)));
  assign y10 = (((b3?p4:a4)-(p1?p2:p5))?((b4?p5:p5)?(b2>=p9):(p7<<<p3)):{(~^(~|p3)),(a0>a2)});
  assign y11 = {(-{a0}),{b5,b1,a2},{a0,b2,a4}};
  assign y12 = (~|(~|{p10,p13}));
  assign y13 = {4{p16}};
  assign y14 = (p14?b3:b3);
  assign y15 = (~&((p9?p17:p15)));
  assign y16 = ((!((-3'sd0)?(5'd3):(~|b5)))^~((-(-5'sd1))<<(p11?p2:a4)));
  assign y17 = (($signed(((p8&p12)<<<$signed(p8)))));
endmodule
