module expression_00244(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(!{(4'sd4),(-4'sd4),(4'd10)}),{(~&(2'd1))}}^~(~^(+((~(-3'sd1))>((-4'sd2)>=(5'd21))))));
  localparam [4:0] p1 = ((|(3'd6))>>>(+(3'd0)));
  localparam [5:0] p2 = ((((3'sd3)|(2'd1))?((4'd8)&&(2'd1)):((3'd4)|(4'd2)))&(((-3'sd2)!==(5'd26))>={(3'd1),(3'd4)}));
  localparam signed [3:0] p3 = ((2'sd0)+(-3'sd1));
  localparam signed [4:0] p4 = {{(5'sd12)},(|(-2'sd1)),{(5'd26)}};
  localparam signed [5:0] p5 = (((3'd7)>=(5'd24))>>{(2'sd0),(3'sd3),(3'd6)});
  localparam [3:0] p6 = (+(^(-{1{{4{(5'sd1)}}}})));
  localparam [4:0] p7 = (2'sd1);
  localparam [5:0] p8 = (((2'sd0)&(2'd1))<<<((-2'sd0)>>(2'd2)));
  localparam signed [3:0] p9 = {2{(|{(((5'sd8)+(3'sd1))|(2'd0))})}};
  localparam signed [4:0] p10 = ((2'sd1)?(4'd15):{4{(-2'sd0)}});
  localparam signed [5:0] p11 = ((((3'sd3)>(4'sd0))<<((5'd12)<=(3'd7)))<=({1{(4'sd1)}}>>>{1{(2'd1)}}));
  localparam [3:0] p12 = (+((4'sd0)?(3'd6):(4'd11)));
  localparam [4:0] p13 = ((-5'sd12)+(5'sd3));
  localparam [5:0] p14 = ((((2'sd0)||(2'd0))<=((2'sd1)>>>(5'd4)))!=((4'd2 * (2'd0))===((5'd1)|(-2'sd1))));
  localparam signed [3:0] p15 = ((2'sd1)^~(3'd0));
  localparam signed [4:0] p16 = {{{(-4'sd6),(2'd0),(4'sd6)}},((4'd8)&&(2'd0))};
  localparam signed [5:0] p17 = {2{(3'd6)}};

  assign y0 = (!(~&((^{4{a4}})!=={(5'd2 * a2),{2{b5}},{3{a2}}})));
  assign y1 = (-((-{(+(~^p15))})?{(a2&p12),{b5},(p4||p13)}:(~{p6,a3,b2})));
  assign y2 = ((^(&{{a4,b1},(p16?b5:p12),{a1}}))<<<(~((a1===a1)^~(a1?b4:a2))));
  assign y3 = (+(p2?p9:p15));
  assign y4 = ((~(a0?a5:a2))?(+(a0?b5:b4)):(!(^(+(&b2)))));
  assign y5 = (({1{(a4<b2)}}!==(b5^~b4))==({4{p11}}<<$signed((p13))));
  assign y6 = ({2{(~^a1)}}|((4'sd2)!=(~p13)));
  assign y7 = (~(~^((-{p2,p14,b2})<<<$signed((-a1)))));
  assign y8 = {2{{{3{b3}},(4'd12)}}};
  assign y9 = (~&($signed({(~^(b5|a4)),(~^(p6>a1)),((p15|p3))})^(((a0!==b3)<<<(a2<<<p7))<=((~^a2)<=(p9<=p12)))));
  assign y10 = (((+(b3===a1))-(^(+p15)))-((p17==a1)-(^(p15>=a3))));
  assign y11 = (2'd2);
  assign y12 = (~&(~^(&(|((-(~|(p6-p11)))?(4'd14):(-5'sd6))))));
  assign y13 = ((!{1{{3{(b1?a4:a2)}}}})^~((a2>>>b0)?(b4?a4:b4):{1{(b0!=b4)}}));
  assign y14 = (-(({p10,b5,p13}^~(a0!==b4))|((^a3)>>>(~&a0))));
  assign y15 = $unsigned((-3'sd3));
  assign y16 = ({(b5?a0:a0),(+b2)});
  assign y17 = (~^(-((6'd2 * (~(a2?a2:p1)))?{2{(b5>b4)}}:((-b2)^(a2^b3)))));
endmodule
