module expression_00908(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^{{(5'sd5),(5'd16)}});
  localparam [4:0] p1 = ((-4'sd2)?(4'd12):((4'd6)==(5'sd3)));
  localparam [5:0] p2 = (5'd2 * (3'd6));
  localparam signed [3:0] p3 = {({{(2'sd1),(3'd1)},((2'd2)>=(4'd13)),{(3'sd2),(5'sd11),(2'sd0)}}||(4'sd2))};
  localparam signed [4:0] p4 = {2{(+{3{(5'd3)}})}};
  localparam signed [5:0] p5 = ({((4'd7)?(3'd3):(-5'sd1)),((-5'sd2)?(-4'sd0):(5'd2))}=={4{{3{(5'sd14)}}}});
  localparam [3:0] p6 = (-4'sd3);
  localparam [4:0] p7 = {3{(3'sd0)}};
  localparam [5:0] p8 = (-5'sd11);
  localparam signed [3:0] p9 = (&(!(~|({(4'sd3),(5'sd15),(5'sd9)}&{(4'd14),(2'sd1)}))));
  localparam signed [4:0] p10 = (2'd2);
  localparam signed [5:0] p11 = (4'd6);
  localparam [3:0] p12 = ((&((4'sd4)?(5'd12):(5'd4)))?(+({2{(5'd14)}}&&(-5'sd13))):(((-3'sd0)?(2'd1):(3'd4))===(~&(-3'sd0))));
  localparam [4:0] p13 = ({2{(!(3'sd2))}}&(~|((^(2'd2))!={1{(5'sd8)}})));
  localparam [5:0] p14 = {3{{3{(2'sd1)}}}};
  localparam signed [3:0] p15 = (5'sd3);
  localparam signed [4:0] p16 = ({(4'd1)}||(|(4'sd0)));
  localparam signed [5:0] p17 = ((((2'd3)==(4'd13))<<((3'd5)>>>(-4'sd5)))<=(~&(+(~&((5'd24)!==(3'sd1))))));

  assign y0 = (~p12);
  assign y1 = (+{{{3{{4{p8}}}}},({p1,p15}?(p0?p5:p2):(p5?p4:p0)),({4{p4}}?{3{p14}}:(~^p6))});
  assign y2 = (~|{1{(&((-4'sd5)))}});
  assign y3 = {(p13<<<a2),(b0!=a2)};
  assign y4 = (b2?a2:a2);
  assign y5 = ({3{(a0==a2)}}&((a2&&p14)>(b4!==b1)));
  assign y6 = (^{(!(&(!(p17^a5))))});
  assign y7 = ((-3'sd0)?(-4'sd3):(~(a5?p11:a1)));
  assign y8 = (5'd26);
  assign y9 = ((~|{4{b3}})|((b5<<<b5)||(p10<=a0)));
  assign y10 = {{a5},(p13-a1),(a4<<a3)};
  assign y11 = {3{((a1^~a5)>>{1{b3}})}};
  assign y12 = {1{b4}};
  assign y13 = (4'sd4);
  assign y14 = {(^(p2^p12)),$unsigned((p11?a5:a5))};
  assign y15 = (((p17<=p10)-(a5>p16))-($signed(p14)?(a4!==a3):(p5-p2)));
  assign y16 = (3'd3);
  assign y17 = {{(4'd2)}};
endmodule
