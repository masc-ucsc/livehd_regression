module expression_00666(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(4'd10)}};
  localparam [4:0] p1 = (({(3'd3),(4'sd0)}?(-(-4'sd0)):((2'd3)?(5'd7):(2'sd1)))===(~({(5'd1),(5'sd10)}^~((4'd9)?(-2'sd1):(-4'sd3)))));
  localparam [5:0] p2 = (|{4{{1{(~^{3{(3'sd2)}})}}}});
  localparam signed [3:0] p3 = ((5'd14)>>>{(-(4'd13)),(|(-(4'd10)))});
  localparam signed [4:0] p4 = (~{4{(-3'sd1)}});
  localparam signed [5:0] p5 = ((|(^((-2'sd0)/(5'sd1))))<<(((-2'sd1)-(-4'sd6))==(~&(5'sd5))));
  localparam [3:0] p6 = ({4{(2'd3)}}^(^(((5'd24)>>(3'd1))||(~(-4'sd7)))));
  localparam [4:0] p7 = (({2{(2'd3)}}?{2{(4'sd5)}}:((4'd7)+(3'd3)))^~(|({1{(2'd0)}}>((5'd5)&&(2'd2)))));
  localparam [5:0] p8 = ((-3'sd3)>=(5'd13));
  localparam signed [3:0] p9 = ((5'sd4)?{{3{(-5'sd6)}}}:((-2'sd1)?(2'sd0):(-4'sd0)));
  localparam signed [4:0] p10 = (((2'sd1)?(4'd0):(2'sd1))?((5'sd10)?(5'sd12):(2'd2)):(((5'd30)?(2'd2):(4'd3))|((-2'sd1)>(3'd5))));
  localparam signed [5:0] p11 = (-((4'sd0)<<<(2'd1)));
  localparam [3:0] p12 = ((((-4'sd1)^~(-5'sd6))-((4'd2)?(-3'sd0):(5'd23)))|(5'd2 * ((4'd8)?(3'd5):(3'd6))));
  localparam [4:0] p13 = (((^(3'd3))<={(4'd4)})-((-5'sd10)?(5'd24):(4'd13)));
  localparam [5:0] p14 = (((3'sd0)&&(5'd8))|((3'd7)?(-3'sd3):(5'd24)));
  localparam signed [3:0] p15 = ((|(-(!(-(^((2'd1)?(-5'sd10):(-3'sd2)))))))&&((~|(~&(-5'sd0)))/(-5'sd2)));
  localparam signed [4:0] p16 = ((4'd12)-(2'd1));
  localparam signed [5:0] p17 = ((-2'sd0)>>>{3{((5'sd1)^~(4'd3))}});

  assign y0 = ((~^(p16?p12:p6))?(p6<<<p9):(~|{p3,a0}));
  assign y1 = ((~&{(+(3'd5)),(b3>>>p6)})<<<((a0<<p16)?(b0===a4):(b1?b2:b4)));
  assign y2 = (-((((((b5-b4)>=$unsigned((~^b0))))))));
  assign y3 = {{1{{4{p2}}}},{{1{{p9,b5}}},{p9,p4,p7}},{{b2,p4,b2},{2{p15}}}};
  assign y4 = ((6'd2 * (p6>>p1))+((^{4{p1}})&&(|(4'd2 * b1))));
  assign y5 = {({{b3},(&a4)}&&{(~b5),(6'd2 * p8),{b0,a1}})};
  assign y6 = ((b0<<<a4)!=(a2==a5));
  assign y7 = (3'd7);
  assign y8 = ((-{4{(a0?a1:a1)}})?(!((a2?a0:b3)-(p7-p17))):($signed({2{a4}})<<<{3{a3}}));
  assign y9 = (b5===a0);
  assign y10 = {3{(~|p13)}};
  assign y11 = (({p3,p12}<<(~|(+p9)))>>{((p2-p11)+(~|p6))});
  assign y12 = (p12>=b4);
  assign y13 = (3'sd2);
  assign y14 = ((2'sd1)<=(~^p4));
  assign y15 = ((((b0>=b5)>(2'd0))==((|a5)||(a3==a4)))!==(((~a5)||(+a0))^~(3'd0)));
  assign y16 = {4{p13}};
  assign y17 = ({(a0^b5)}===(~(a5<b5)));
endmodule
