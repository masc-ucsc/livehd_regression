module expression_00406(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&{2{(-2'sd0)}});
  localparam [4:0] p1 = (+(((3'd5)||(4'd5))==((3'd6)+(2'd0))));
  localparam [5:0] p2 = {4{(5'sd2)}};
  localparam signed [3:0] p3 = (&(2'd2));
  localparam signed [4:0] p4 = ((~(+(3'd5)))%(2'd1));
  localparam signed [5:0] p5 = (!(-(-(-({2{(^(&(2'd0)))}}>(|((&(4'sd5))==((5'sd12)<<(3'd5)))))))));
  localparam [3:0] p6 = (&(~((~{1{(4'd15)}})?(~|{3{(3'sd1)}}):{4{(3'sd1)}})));
  localparam [4:0] p7 = ({(4'd10),(5'd14)}?((5'd0)===(4'd15)):((3'sd2)<=(4'd1)));
  localparam [5:0] p8 = (((3'd6)==(3'd4))<=(~|((2'd3)>=(-2'sd1))));
  localparam signed [3:0] p9 = (&{4{((4'd2)?(5'sd5):(3'sd3))}});
  localparam signed [4:0] p10 = ({3{(4'd3)}}?((4'd10)>(3'sd2)):((3'd2)?(2'd2):(3'sd0)));
  localparam signed [5:0] p11 = {((2'd2)>=(4'd13)),(-(|(2'sd1))),(~|((5'd4)&&(2'd0)))};
  localparam [3:0] p12 = {(((4'sd1)?(-2'sd1):(5'd30))&&(~^(~^(4'd12))))};
  localparam [4:0] p13 = (((~{3{(-2'sd0)}})>(~(~&(4'd14))))^{3{(~^(5'd22))}});
  localparam [5:0] p14 = (((2'd1)?(2'd1):(4'sd3))?(-4'sd7):{1{(2'sd1)}});
  localparam signed [3:0] p15 = (~|(~&((!(2'd0))=={(-2'sd1)})));
  localparam signed [4:0] p16 = {{(^{(5'sd4),(2'd1)}),(~&(~((3'd5)?(3'sd2):(5'd13))))},{{(((3'sd0)?(-5'sd9):(4'sd5))?{(2'd2),(3'd6)}:{(4'sd2),(2'sd0)})}}};
  localparam signed [5:0] p17 = (((2'd1)?(2'd0):(3'sd1))?((5'd2)&&(5'd15)):((5'sd2)?(-3'sd0):(3'd7)));

  assign y0 = (({1{((a2&b0)&{2{b1}})}}<((b0<b0)<<<{3{p7}}))>(((p5&&p6)<<{1{p10}})==((b3<<b1)!==(4'd2 * a1))));
  assign y1 = {$signed($unsigned({{3{p12}},{{3{p14}}}}))};
  assign y2 = (^(~|(-((a5===b5)?(b2<<<b2):(b1>>p8)))));
  assign y3 = (a0?p12:a2);
  assign y4 = (3'sd0);
  assign y5 = ((b4%p0)?(b1+p12):(b1?b5:p0));
  assign y6 = ({2{(b5?p4:b2)}}?((^p16)?(2'd3):(3'sd0)):(~|$signed((-(b4)))));
  assign y7 = ((p1!=p2)>>>(b1===b4));
  assign y8 = (5'd28);
  assign y9 = (b1&&a4);
  assign y10 = (~|(((b0)<<<(a5||a4))&&(~^(5'sd14))));
  assign y11 = {3{p7}};
  assign y12 = $unsigned({{3{{2{p3}}}}});
  assign y13 = ((2'sd1));
  assign y14 = $unsigned((^(&((^(p3?p6:p16))<<(4'd14)))));
  assign y15 = (5'd0);
  assign y16 = {(((a1?p10:p7)<<<(^a0))?(&{p4,b1,p7}):((b1?p14:b3)+(a0?a2:p12)))};
  assign y17 = ({p0,b4,a5}>=(a5<<p14));
endmodule
