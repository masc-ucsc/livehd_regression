module expression_00050(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(~|(!(((2'd3)>=(5'd22))<{(3'd5),(5'd23),(2'sd1)})))};
  localparam [4:0] p1 = {(^{(~((4'd10)?(5'sd0):(-2'sd0)))}),(((4'd12)!==(-5'sd9))?((2'd3)&&(2'sd1)):{(2'd1)})};
  localparam [5:0] p2 = (|(-{1{{(+{{(3'sd1),(5'sd13),(3'd3)},(!(4'sd2))})}}}));
  localparam signed [3:0] p3 = ((~|(-2'sd0))?{(5'sd0),(5'sd4),(5'sd10)}:{(-3'sd0)});
  localparam signed [4:0] p4 = {(|((+{(-2'sd1),(-4'sd7),(-4'sd0)})<<{((3'd6)?(-3'sd1):(3'd6)),((-4'sd6)?(-2'sd1):(4'sd5)),((4'd12)^~(4'sd2))}))};
  localparam signed [5:0] p5 = (^(5'sd13));
  localparam [3:0] p6 = ((^(5'd6))*(-(5'sd2)));
  localparam [4:0] p7 = {4{(~(-5'sd0))}};
  localparam [5:0] p8 = (((4'sd0)?(-3'sd3):(4'd3))?{4{(-4'sd0)}}:{3{(-3'sd0)}});
  localparam signed [3:0] p9 = ((((2'd1)?(3'd5):(-3'sd2))<=((2'sd1)?(-4'sd3):(-2'sd1)))<(((4'd3)?(5'sd7):(4'd7))?((-5'sd0)>=(3'sd3)):{(-4'sd7),(4'd13)}));
  localparam signed [4:0] p10 = (-(~^(&(~|(((2'd0)?(-4'sd1):(3'd4))?((5'sd15)?(2'sd0):(-4'sd0)):((-3'sd2)?(2'd1):(2'sd0)))))));
  localparam signed [5:0] p11 = ({1{(((5'd31)?(4'd8):(-5'sd3))!=={2{(-4'sd1)}})}}?((^(-4'sd0))<<((-2'sd1)?(4'd0):(2'sd1))):(((-4'sd0)+(3'd6))?((4'd8)?(-3'sd1):(5'd5)):((-4'sd2)^(5'd0))));
  localparam [3:0] p12 = ((5'sd1)?(3'sd1):(-2'sd1));
  localparam [4:0] p13 = (5'd15);
  localparam [5:0] p14 = {{4{(4'd1)}},{(3'sd3),(-4'sd1)},{4{(2'sd1)}}};
  localparam signed [3:0] p15 = ((((-3'sd0)>(2'sd0))>{4{(-4'sd5)}})+(~(~&(~|(^{1{(-4'sd6)}})))));
  localparam signed [4:0] p16 = (((6'd2 * (4'd10))<((4'sd5)<<(3'd6)))>(~(((-4'sd3)>>(4'd15))<=((3'd6)<=(2'd3)))));
  localparam signed [5:0] p17 = (-5'sd13);

  assign y0 = (4'd0);
  assign y1 = (p17?a3:b3);
  assign y2 = (~$signed((~|{{b5,a2,p17},(|({p6})),({p15}|$signed(b3))})));
  assign y3 = (b2?a1:p1);
  assign y4 = (!(-5'sd7));
  assign y5 = (-2'sd0);
  assign y6 = (((b5>>>b1))/b1);
  assign y7 = {3{((-5'sd14))}};
  assign y8 = (~(((-p12)&(~|p11))<(~|(p12-b5))));
  assign y9 = {4{(4'sd5)}};
  assign y10 = (~|(-(~|(+(~|((+($signed(b2)!==(~&a1)))|(~|(~^(4'd2 * p8)))))))));
  assign y11 = {1{({2{((b3>>a2)<<<(~&a1))}})}};
  assign y12 = (((a5+a0)%a0)<<<(~^((+b4)^~(~&a0))));
  assign y13 = $unsigned(((({3{p0}}|(2'd2))||(-5'sd11))&&{4{(a4<<<p0)}}));
  assign y14 = (&(+{2{(!(+{3{{4{p15}}}}))}}));
  assign y15 = (-((&(~|p0))));
  assign y16 = (((~|b5)||{a0})>$signed({b0,p12,b3}));
  assign y17 = (((b5?p17:p17)?(p3?p16:b0):(p14>=p17))?((b1?p10:p7)/p17):((p16?p7:p0)<(p10?p6:p9)));
endmodule
