module expression_00484(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd22)<=(3'd3));
  localparam [4:0] p1 = {4{(&(~|{4{(2'd3)}}))}};
  localparam [5:0] p2 = {1{((+{2{(-(2'd1))}})>>>{(-(4'd3)),(~|(-4'sd2)),{(5'd7)}})}};
  localparam signed [3:0] p3 = (5'd2 * ((5'd22)&(2'd0)));
  localparam signed [4:0] p4 = ((((3'd1)^(4'd1))&((2'sd1)||(5'd12)))<=(((-2'sd0)^(3'd2))||((4'sd3)<<(5'sd8))));
  localparam signed [5:0] p5 = {1{(~|((-5'sd10)||(3'd6)))}};
  localparam [3:0] p6 = {3{(4'd1)}};
  localparam [4:0] p7 = (^(4'd3));
  localparam [5:0] p8 = {3{{1{(|((2'sd1)!==(4'd8)))}}}};
  localparam signed [3:0] p9 = ({1{((-4'sd4)||(4'd2))}}|(-(+(3'd1))));
  localparam signed [4:0] p10 = {2{{2{((5'd13)?(-2'sd1):(4'd4))}}}};
  localparam signed [5:0] p11 = (3'd6);
  localparam [3:0] p12 = (&(-4'sd2));
  localparam [4:0] p13 = ((^(-5'sd8))>>(&(!(-4'sd1))));
  localparam [5:0] p14 = ({4{(|(2'sd0))}}===(((3'sd3)?(-5'sd2):(3'd5))?(^(5'd1)):((4'd13)|(5'd6))));
  localparam signed [3:0] p15 = (4'd9);
  localparam signed [4:0] p16 = {1{((((2'd2)-(-2'sd1))?((2'sd1)<=(2'd3)):((2'd2)?(2'sd0):(3'd5)))!=={2{{1{{2{(4'sd7)}}}}}})}};
  localparam signed [5:0] p17 = {4{((2'sd0)?(5'd6):(5'sd4))}};

  assign y0 = (p10);
  assign y1 = (3'sd2);
  assign y2 = ({4{{b5,b0}}}^~(4'd2 * {b0,p8,a1}));
  assign y3 = {(5'd30),(6'd2 * (p0^b0)),(4'd8)};
  assign y4 = (((p16?p2:b0)^(2'sd1))<<((a2>>>b1)>>>(b4%p2)));
  assign y5 = (p11&p10);
  assign y6 = (($unsigned((~p7))<(a5*b3))<(~^($unsigned((a0!==b2))>((|b3)))));
  assign y7 = {1{{3{(&{4{b4}})}}}};
  assign y8 = {(~(~^(~|{1{b5}}))),(~^(~(a4!=a2))),((b3!=b1)-{b0,p2})};
  assign y9 = ((-2'sd0));
  assign y10 = (-3'sd3);
  assign y11 = {3{{2{p13}}}};
  assign y12 = ((4'd7)<<(~^a3));
  assign y13 = (-{2{{1{(+(-2'sd1))}}}});
  assign y14 = {p17};
  assign y15 = ((~|(2'd2)));
  assign y16 = ({3{(b2>>b4)}}==(((~^b0)||(+p8))+{4{b4}}));
  assign y17 = ((b4<<<b5)*(p10>=b1));
endmodule
