module expression_00308(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{((3'd1)+(4'sd2))}};
  localparam [4:0] p1 = (((3'd2)^~(4'd10))+{(5'd24),(3'd0),(-3'sd1)});
  localparam [5:0] p2 = (-((~|((4'd6)&(5'd14)))==(|(!((2'd1)?(3'd6):(3'd3))))));
  localparam signed [3:0] p3 = (|((3'sd0)<=(3'd5)));
  localparam signed [4:0] p4 = (((5'd9)<<(2'sd1))<((5'sd0)<(2'd0)));
  localparam signed [5:0] p5 = (^(5'sd2));
  localparam [3:0] p6 = {2{(((4'd12)>>(5'd3))&((2'sd1)&&(3'sd1)))}};
  localparam [4:0] p7 = (((3'd4)|(4'd8))>((5'sd3)+(3'sd1)));
  localparam [5:0] p8 = (((~&((-2'sd0)|(2'sd1)))>{(5'sd9),(2'd3)})>>>{1{(!({(-5'sd6),(-5'sd5),(3'd0)}==((5'd9)>=(-3'sd3))))}});
  localparam signed [3:0] p9 = (((3'd3)>>>((3'd0)||(-4'sd4)))?(((-5'sd7)>=(4'd9))===((4'sd5)|(3'sd2))):((-(-5'sd13))&(~(4'd9))));
  localparam signed [4:0] p10 = ((2'sd1)^(-3'sd1));
  localparam signed [5:0] p11 = (4'd2 * (&((2'd1)|(2'd3))));
  localparam [3:0] p12 = (((-3'sd0)?(5'd16):(-4'sd3))<<<((5'd24)?(5'd4):(-4'sd6)));
  localparam [4:0] p13 = ((4'd0)?(5'd28):(3'sd1));
  localparam [5:0] p14 = ({(~^{1{((-4'sd4)?(5'd31):(5'sd7))}})}?((+(3'sd2))?{(5'd13),(2'sd1),(-3'sd2)}:((-3'sd2)?(4'd2):(3'sd1))):(2'd3));
  localparam signed [3:0] p15 = (~|(5'd23));
  localparam signed [4:0] p16 = ((4'd2 * {1{((5'd23)>(3'd0))}})>{3{{3{(-3'sd3)}}}});
  localparam signed [5:0] p17 = (2'sd1);

  assign y0 = (&(~^(^{{p10,p8,p0}})));
  assign y1 = (3'd2);
  assign y2 = {3{{1{(2'd1)}}}};
  assign y3 = (p16==p10);
  assign y4 = ((~&(a2<=p12))<=((a4==b1)));
  assign y5 = (((~^(b0<p8))-{1{(b1>b1)}})<((p8&&a1)>=$signed({1{b5}})));
  assign y6 = ($signed(($unsigned(b4)>>(b4|b0)))>=((a4)&(a1<=b3)));
  assign y7 = (p1<<<b0);
  assign y8 = {$unsigned({({p14,a0}),(+$signed(a5))}),{$signed((b5===b4)),{1{(b1<a3)}}},{4{(b4>>>b4)}}};
  assign y9 = $signed($unsigned((&(~^(+((b3>=p4)?(b2?a4:b0):(^a1)))))));
  assign y10 = (~((~&((p8?p11:p14)>>(p10?p7:p16)))?((a0?a0:b5)!==(b5===b0)):(|(p0?p7:p1))));
  assign y11 = (~^$unsigned({(2'd1),$signed({(+(!$signed(p0)))})}));
  assign y12 = (a5?a3:b0);
  assign y13 = {3{(({3{b5}})^(^(a3&&p16)))}};
  assign y14 = ({p13,b0,b3}<(b1?a4:a1));
  assign y15 = {2{(~&p9)}};
  assign y16 = (2'sd0);
  assign y17 = ((5'd19)>>>((4'd2 * p6)<<<(p9?p13:p9)));
endmodule
