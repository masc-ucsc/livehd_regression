module expression_00136(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(4'd1)}};
  localparam [4:0] p1 = (-3'sd3);
  localparam [5:0] p2 = (^(~&{{{((~(5'd3))&&((-2'sd1)===(3'd0))),(~^({(3'd7)}|(~&(3'd2))))}}}));
  localparam signed [3:0] p3 = ((5'd31)-(5'sd2));
  localparam signed [4:0] p4 = ((3'd1)||({(2'sd0),(3'd3)}^~((3'd2)|(3'd6))));
  localparam signed [5:0] p5 = (((4'd12)+(2'd3))||((4'd13)&&(4'd2)));
  localparam [3:0] p6 = ((((4'd12)|((4'sd4)!==(2'sd0)))<{((5'd9)<(-2'sd1)),((5'd18)?(-5'sd15):(4'sd7))})>>(~|(!({1{((3'd2)||(-5'sd5))}}||((-2'sd0)?(2'd1):(-5'sd4))))));
  localparam [4:0] p7 = ((&(&(3'd3)))*(-(-(-2'sd0))));
  localparam [5:0] p8 = {((~|{(4'd14),(3'd2)})^((3'd0)>=(2'd3)))};
  localparam signed [3:0] p9 = (3'sd1);
  localparam signed [4:0] p10 = ((((4'd1)?(-5'sd11):(2'd0))<={(-4'sd7),(4'd3)})==(-(!((3'd4)?(5'sd15):(2'sd0)))));
  localparam signed [5:0] p11 = (((|(4'sd6))?((3'sd1)/(3'd7)):((5'sd9)!=(4'sd3)))<<((&(5'd1))?(&(-3'sd2)):((-2'sd1)?(2'd2):(4'd9))));
  localparam [3:0] p12 = ((4'd4)<(4'd14));
  localparam [4:0] p13 = (2'd2);
  localparam [5:0] p14 = (3'd7);
  localparam signed [3:0] p15 = (5'd1);
  localparam signed [4:0] p16 = (4'd5);
  localparam signed [5:0] p17 = (2'd1);

  assign y0 = ({p13,p8}!={(3'd5)});
  assign y1 = (($signed(((p10&&p2)<<(+p1)))-(3'd3))&(((5'd0)&(~^(p1%p16)))));
  assign y2 = {3{({1{(p2)}}<<<((p8>p8)))}};
  assign y3 = $unsigned({3{p10}});
  assign y4 = {3{(&{a3,p0,a0})}};
  assign y5 = $signed(($signed(((!b4)^(a1<<<a4)))<=((p5>a0)>>{4{a1}})));
  assign y6 = ({$signed((~(b0-a0)))});
  assign y7 = (4'd12);
  assign y8 = {2{({4{b3}}?(+{2{p11}}):(~^{4{b5}}))}};
  assign y9 = (&{1{((~{1{(2'd3)}})===(4'd13))}});
  assign y10 = (((a5&&a4)+{a3})!==(5'sd13));
  assign y11 = (((-(~|(4'd2 * a1)))===(~&(+(b0>a0))))>=(2'd0));
  assign y12 = (+(a3+a4));
  assign y13 = ((~|{2{{2{{4{p7}}}}}})||(2'd0));
  assign y14 = ((2'sd0)?((4'd9)?(4'd3):{b3,a0,a3}):((a5?a5:a0)?{a1}:{a5}));
  assign y15 = ({1{b0}}?(a4+a0):(p10?a4:b4));
  assign y16 = (~(^(((-a2)<<<{1{b2}})<={2{(a0<<b4)}})));
  assign y17 = ((((a3||b3)!=(b5===b5))!==((b1==a1)<<(b2^~a5)))>(((b2*b3)*(p13&&b0))^~((a3<<a5)===(b2<=b5))));
endmodule
