module expression_00654(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'sd9)^((4'd1)|(3'd4)));
  localparam [4:0] p1 = (-(-((+(|(2'sd1)))%(-4'sd3))));
  localparam [5:0] p2 = ((5'd20)-(5'd5));
  localparam signed [3:0] p3 = {(((-5'sd7)&&(2'd3))+((4'd12)+(3'd0))),({1{(2'd3)}}!=((2'd2)&&(4'sd6))),{((3'sd3)^(2'sd0))}};
  localparam signed [4:0] p4 = (((-2'sd0)>>(5'd16))>(~&((-3'sd0)-(4'sd0))));
  localparam signed [5:0] p5 = (((5'd0)?(5'd25):(3'd0))?((-3'sd0)!=(-2'sd0)):((3'd2)?(4'sd0):(3'sd3)));
  localparam [3:0] p6 = ((~(((5'd17)?(5'd16):(3'd3))>((4'sd2)+(3'sd2))))===(^(~{(3'd1)})));
  localparam [4:0] p7 = (^{((5'sd2)!=(3'd6)),((5'sd9)>(5'sd5)),(4'd1)});
  localparam [5:0] p8 = (!(&(&(+(&(&(~|(4'd0))))))));
  localparam signed [3:0] p9 = (((3'd4)?(4'd5):(4'd5))?(~&(5'd6)):(&(4'd7)));
  localparam signed [4:0] p10 = {2{{1{{2{(3'd0)}}}}}};
  localparam signed [5:0] p11 = (!(+(~(~&((&((~(-2'sd1))+((2'd3)!=(3'd6))))<<(~|(&(4'd2 * (3'd4)))))))));
  localparam [3:0] p12 = (^{(~^{(-3'sd0),(5'd25)}),{(2'd0),(4'sd3),(2'sd1)},(~&{(-5'sd14)})});
  localparam [4:0] p13 = (~^(((2'd2)?(5'd10):(-2'sd1))?(~|((2'd2)?(5'd18):(5'd15))):((-4'sd7)?(-4'sd3):(5'd21))));
  localparam [5:0] p14 = (((4'sd4)===(5'd2))-((-3'sd1)>>(4'd3)));
  localparam signed [3:0] p15 = (^(&(2'd0)));
  localparam signed [4:0] p16 = ((5'd6)<<(((3'd3)*(5'sd11))<<((-5'sd6)!=(5'sd5))));
  localparam signed [5:0] p17 = ((~|(-5'sd4))&&{4{(4'sd7)}});

  assign y0 = {2{(~^(b4<=a0))}};
  assign y1 = (4'd2 * (p12^~b0));
  assign y2 = (((4'd2 * (a2>a2))<={b1,b0,a2})^{({{b5,b0,b2}}<{(a2^b2),(a1>>>a0)})});
  assign y3 = (({(a5==b5),{p0}}!=(!{(b3>>a4)}))>=(((^p11)==(!b1))>>{(a0==b0)}));
  assign y4 = {2{(^((-4'sd2)?{1{b4}}:(|b2)))}};
  assign y5 = ((~&{2{{2{p16}}}}));
  assign y6 = (&{3{{2{p11}}}});
  assign y7 = {4{(p17?p7:p6)}};
  assign y8 = (((4'sd4)));
  assign y9 = (((a2*b4)^(a1?a2:b3))>((b2?b3:b5)<=(a2*b4)));
  assign y10 = {(5'd29),((2'd0)&(&{1{(2'd0)}}))};
  assign y11 = {p14};
  assign y12 = (~((a2>a5)!==(a3+b3)));
  assign y13 = {3{(|{3{(p15&p1)}})}};
  assign y14 = {2{{p11,p7,b2}}};
  assign y15 = ((|(&(p8+a3)))?(^(~^(~|p12))):((b3&b0)*(p9%p17)));
  assign y16 = (~^(-(~|(^(^$signed($unsigned((|((~^(!$signed($signed($unsigned((-(^p0))))))))))))))));
  assign y17 = ((-{p7,p17,a4})<<{p5,b0,b3});
endmodule
