module expression_00472(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{((5'd2)!==(2'd2))}};
  localparam [4:0] p1 = {((-2'sd1)&&(-5'sd15))};
  localparam [5:0] p2 = ((2'd1)<<<(5'd20));
  localparam signed [3:0] p3 = {4{((~|(3'd2))>=((-3'sd1)&&(2'd1)))}};
  localparam signed [4:0] p4 = ((~((|(-4'sd0))>((3'sd2)==(3'sd1))))<(((5'sd6)>>(2'd1))>>>(|(^(3'd6)))));
  localparam signed [5:0] p5 = (-5'sd13);
  localparam [3:0] p6 = {(~^(-4'sd1)),{(-5'sd15)},(^(4'd0))};
  localparam [4:0] p7 = ((-(-{2{(-4'sd5)}}))>(|((4'd3)<<(4'sd4))));
  localparam [5:0] p8 = (&(((5'sd1)<<(5'sd6))<=((4'd6)!=(5'sd1))));
  localparam signed [3:0] p9 = {2{(-(2'd2))}};
  localparam signed [4:0] p10 = (&(&((4'd14)?(-2'sd1):(3'sd3))));
  localparam signed [5:0] p11 = {(~&((-3'sd2)-(-4'sd6))),{(3'd5),(5'd9)},((2'd3)>>>(2'sd0))};
  localparam [3:0] p12 = {(((5'd27)?(5'd11):(2'd0))?(^((5'd2)?(2'sd0):(4'd10))):((2'sd1)?(4'd2):(5'sd3)))};
  localparam [4:0] p13 = ({1{((-3'sd1)-(4'sd6))}}-{(-5'sd14),(-2'sd1),(4'd2)});
  localparam [5:0] p14 = {(-(~&(4'sd1))),{((5'd8)>>>(-5'sd13))},(^((-3'sd0)?(5'd6):(5'd11)))};
  localparam signed [3:0] p15 = (2'd1);
  localparam signed [4:0] p16 = {1{(4'sd1)}};
  localparam signed [5:0] p17 = (((-2'sd0)<=(2'd1))===(4'd0));

  assign y0 = (((^(a0+p3)))?((+b0)*$unsigned(b2)):(p15?b2:p7));
  assign y1 = ((4'd2 * (|(b1^~a0)))===({4{b1}}>>{4{a4}}));
  assign y2 = ((-(b3^~a5))?(~&(4'd0)):((b2&b3)||(~|p17)));
  assign y3 = (^(-5'sd7));
  assign y4 = (|((&(p12|p12))==(p0?p9:p16)));
  assign y5 = {(&{4{(~&(!b1))}})};
  assign y6 = $signed((-4'sd3));
  assign y7 = (({a2,b0,a0}>>{a5,a1})?{{b4,a1,b1},(a5?a5:a5)}:{{2{(b3^b0)}}});
  assign y8 = (5'sd4);
  assign y9 = {({3{(~{1{a1}})}}^~{{{2{b4}},(6'd2 * p0)},{2{(p12?a1:p11)}}})};
  assign y10 = {(b1||p8)};
  assign y11 = ({2{(a1>b2)}}?({p14}?{p15,b4}:$unsigned(p14)):{(4'd7),(a0?p15:p1)});
  assign y12 = {1{{3{((p13?p13:a1)<=$signed((a0?b4:a1)))}}}};
  assign y13 = (-5'sd8);
  assign y14 = ({3{(p10<<<p4)}}>>>({1{(p8^b5)}}!=(p1>>>p10)));
  assign y15 = (((&(4'd3))>>(b3?p12:a4))<=((5'd2 * a0)^(-4'sd2)));
  assign y16 = {3{p16}};
  assign y17 = ({{1{(a4<<p6)}}}||{1{{{2{b3}},(a4<b2)}}});
endmodule
