module expression_00347(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|{{((-2'sd0)>>(2'd3))},(!(~((2'd3)==(4'sd2)))),{{{(3'd3)}}}});
  localparam [4:0] p1 = (((3'sd2)?(5'sd6):(3'd7))>>((5'd29)>>(3'd1)));
  localparam [5:0] p2 = {(((-4'sd4)<(4'sd7))!==(+(5'sd2))),{(3'd7),((4'd7)?(2'd2):(5'sd0)),(&(3'd6))}};
  localparam signed [3:0] p3 = (2'd2);
  localparam signed [4:0] p4 = ((4'd7)?{1{(4'sd5)}}:((-3'sd1)^~(-2'sd1)));
  localparam signed [5:0] p5 = ({(((-5'sd11)^~(2'd1))^~{(-4'sd4)})}=={{((3'd3)^~(-4'sd7)),((5'd14)||(4'd7))}});
  localparam [3:0] p6 = ((&{1{((-5'sd9)?(5'd15):(-3'sd2))}})+{4{(4'd10)}});
  localparam [4:0] p7 = ((+(&(-2'sd0)))>(((5'd14)<<(4'sd0))<<(&((5'sd0)<=(2'd3)))));
  localparam [5:0] p8 = (5'd2 * (~&((3'd5)<<(2'd2))));
  localparam signed [3:0] p9 = {((5'sd2)?(3'd3):(-5'sd6)),(3'd7),{(4'd0),(2'sd0),(3'd7)}};
  localparam signed [4:0] p10 = ({(4'd1),(2'd2),(2'd3)}|{2{(-3'sd3)}});
  localparam signed [5:0] p11 = (~^((5'd2 * ((2'd2)-(2'd2)))?(((4'd7)-(-4'sd0))&((5'd8)?(5'd7):(4'd12))):((+(4'd5))*(~^(-3'sd1)))));
  localparam [3:0] p12 = (((3'd6)^~(-5'sd1))==(2'sd0));
  localparam [4:0] p13 = {3{(4'd8)}};
  localparam [5:0] p14 = ((~(-3'sd3))^((5'd26)?(-3'sd2):(4'd13)));
  localparam signed [3:0] p15 = {(+(5'sd8)),((5'd1)||(-4'sd5))};
  localparam signed [4:0] p16 = {(4'sd3),(-2'sd1),(5'sd4)};
  localparam signed [5:0] p17 = (({(5'sd10),(5'sd6),(5'd1)}<((3'd3)<<(5'sd10)))||((^((5'd28)!==(5'd7)))<<(4'd4)));

  assign y0 = (((&$unsigned((4'd2)))^(3'd5))===(~|(~|(+((!(-2'sd1))-(a2>=a1))))));
  assign y1 = {4{(-(~&(p11?p4:p1)))}};
  assign y2 = ((a2?b4:b0)/b4);
  assign y3 = ($signed((+($signed($signed(p15))||(^(p12^~b0)))))>>>(({b2,p4}<={a2,p13})<((p5)<{p9})));
  assign y4 = ({((a4?b0:b1))}?(4'd2 * $unsigned(b4)):(a5?a1:a4));
  assign y5 = (&{$signed((~|((~^b0)))),(((a3|a0)))});
  assign y6 = ({1{(a1?a3:a2)}}?((-3'sd2)<<<(a3?a3:a5)):((b0^~a1)>>{3{b5}}));
  assign y7 = ((((p6<p2)<<(p6>=b2))>>>((b5?a5:b1)===(4'd2 * a1)))||(((p13?p3:a3)|(6'd2 * p0))-{1{(p15^~b5)}}));
  assign y8 = ((a5==b3)!==(a0||b1));
  assign y9 = (((+(~&(!p7)))>=((~&p2)^~(+p2)))|{((p12!=p7)!={(~|b5)})});
  assign y10 = ((2'sd1)^~(~&(4'd10)));
  assign y11 = ((~^(~|((a2-b2)>(b3*p11))))-((~&(b2|a4))!==((b0==b3)<<(!a3))));
  assign y12 = {3{((p17?a5:p8)<<<(b3<<b5))}};
  assign y13 = (((b4||b3)?(a5?p7:p12):(p3?a1:p11))?((a3===a5)?(b4?a4:p13):(p3?b4:p9)):((b2?a2:a0)==(p15?b2:a2)));
  assign y14 = ((&{(b5!=p6),{2{b2}},(6'd2 * a1)})-((a3|a5)<($unsigned(b3))));
  assign y15 = (4'd3);
  assign y16 = (~|(p2+p14));
  assign y17 = (|(~(!((+p9)?(!a2):(^p16)))));
endmodule
