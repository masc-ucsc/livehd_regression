module expression_00342(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-4'sd5)?(4'd15):(3'd4))?((2'd2)?(2'd0):(4'd2)):((5'd7)?(2'd0):(4'd13)))?(4'd9):(2'd0));
  localparam [4:0] p1 = (((-3'sd2)!==(2'd1))^~((4'd9)&(4'd14)));
  localparam [5:0] p2 = (~&((~|((-5'sd12)+(2'sd1)))==(!((2'sd1)>=(-5'sd4)))));
  localparam signed [3:0] p3 = ((!((-3'sd3)?(5'sd13):(-2'sd0)))<(((3'd0)?(2'd0):(5'sd8))<={1{(3'd3)}}));
  localparam signed [4:0] p4 = (-((~|((4'd1)===(-3'sd3)))===((-4'sd6)+(3'd3))));
  localparam signed [5:0] p5 = ((~^(+(((3'd4)/(-5'sd1))||((3'd2)===(2'd0)))))<<<(|(+(!((-5'sd1)==(2'sd0))))));
  localparam [3:0] p6 = ({3{{2{(3'd4)}}}}===(((-4'sd3)^(2'd3))+((2'd0)-(4'd0))));
  localparam [4:0] p7 = ({(3'd2),(4'd4)}<=((5'sd11)<=(3'd0)));
  localparam [5:0] p8 = (~&((((4'd5)==(5'd17))+{(5'd13),(5'd3)})?(-{(-4'sd5),(-5'sd1)}):((|(-3'sd3))=={(-3'sd2),(-4'sd3),(3'd5)})));
  localparam signed [3:0] p9 = {{((-3'sd2)<(2'd0))},((2'd1)?(3'sd1):(4'd15)),{1{{(2'd1)}}}};
  localparam signed [4:0] p10 = ((((-2'sd0)||(4'd8))>>>((5'd31)===(5'd31)))!==(5'd2 * ((3'd7)^(3'd0))));
  localparam signed [5:0] p11 = ((&((5'sd10)==(4'd8)))!=(-((2'd1)<=(-3'sd1))));
  localparam [3:0] p12 = (((((3'd6)?(3'sd2):(-5'sd3))<=(~(4'sd5)))!==(((2'sd1)==(3'd5))|((-4'sd6)?(-4'sd4):(5'sd2))))>=((~((-5'sd1)>(2'd0)))?((-4'sd3)^~(2'd2)):((4'd2)>(2'sd0))));
  localparam [4:0] p13 = (((+(&(2'd3)))>>>((5'sd12)<(5'd2)))>>>(((2'd1)>(4'd12))-((-2'sd0)===(3'sd1))));
  localparam [5:0] p14 = ((-(5'd31))+(^(4'sd1)));
  localparam signed [3:0] p15 = ((((2'sd0)?(4'd0):(3'sd1))?((3'sd3)>>(3'd6)):((2'd1)?(3'd2):(-2'sd0)))^{{(|(5'd31)),(~&(5'd23))}});
  localparam signed [4:0] p16 = ((4'd13)==(-4'sd6));
  localparam signed [5:0] p17 = ((-5'sd13)>>>(5'd21));

  assign y0 = ((b2==b4)%a1);
  assign y1 = {4{{2{b4}}}};
  assign y2 = (2'd1);
  assign y3 = ({{4{p2}},(-4'sd3)}<<(2'd0));
  assign y4 = $unsigned((((3'd3)?(5'sd7):(p8?p17:p14))));
  assign y5 = {2{{(~^(~b4)),{(p2?p13:b0)},(~(p2))}}};
  assign y6 = ((6'd2 * $unsigned(p9))?$signed($unsigned((4'd7))):$signed($signed((b3&a2))));
  assign y7 = {{(|{(p3<<a5),{p14,b5},(p5>=p6)}),(((&b3)!=(a0-a2))!==(~&(~&(+{a2,b3,b4}))))}};
  assign y8 = ((a0|a0)<<<(b2===b2));
  assign y9 = $signed({4{$unsigned($signed({b0,p2}))}});
  assign y10 = (((&p8)<=(4'sd7))>(^(p6||p5)));
  assign y11 = {(-5'sd5)};
  assign y12 = ((a3&b4)&&((p7^~b2)));
  assign y13 = $signed((5'd3));
  assign y14 = (&(~|((4'd2 * {b1,b2,b0})?((a4-a2)?(a4?a2:b5):(b1?b0:a5)):{1{{1{(p10?b1:a2)}}}})));
  assign y15 = {(-p14),(4'sd1),(2'd2)};
  assign y16 = (((p14?p4:p15)||(p2&&p5))?(5'd2 * (p0?p7:p13)):(2'd2));
  assign y17 = (~&{2{{4{a1}}}});
endmodule
