module expression_00557(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'd3),(2'd3),(3'd6)};
  localparam [4:0] p1 = (+{{(~((-3'sd0)!=(4'd5))),((-2'sd1)!=(2'd0))},(~^((5'd6)&&(^(2'sd0))))});
  localparam [5:0] p2 = {(5'd2 * {3{(3'd7)}})};
  localparam signed [3:0] p3 = (({3{(-4'sd3)}}<=((3'd3)+(2'd1)))&&{(-3'sd3),(5'sd7),(4'd6)});
  localparam signed [4:0] p4 = (~^(-(~&(((2'd2)?(5'd0):(2'd3))==((-2'sd1)!=(3'd2))))));
  localparam signed [5:0] p5 = (&(5'd30));
  localparam [3:0] p6 = (+(((-4'sd5)?(5'sd1):(4'd12))!=(~&((2'd0)>(-5'sd6)))));
  localparam [4:0] p7 = (((5'sd3)?(-3'sd0):(-2'sd0))?{1{(-3'sd1)}}:((5'd20)?(3'sd1):(-4'sd1)));
  localparam [5:0] p8 = {((^((3'sd1)!=(5'sd0)))>=(3'd4))};
  localparam signed [3:0] p9 = (!(((^(4'd14))>=((4'sd4)^~(4'sd5)))^~(5'sd13)));
  localparam signed [4:0] p10 = (^{1{(+{4{((4'sd4)<<(5'd12))}})}});
  localparam signed [5:0] p11 = ((((-2'sd0)+(3'd6))^~((2'd3)>=(3'd6)))?(((3'd2)===(5'd28))+(~(4'd7))):(3'd5));
  localparam [3:0] p12 = (&((((5'd15)>>(-3'sd3))?((3'sd2)&&(3'sd3)):(5'd2 * (5'd10)))-(((2'd0)?(3'd5):(4'sd4))<<<((3'sd3)>(5'd9)))));
  localparam [4:0] p13 = ((((2'd3)!==(4'd9))?((-2'sd1)?(2'd1):(5'd23)):((-2'sd1)==(5'sd8)))|(6'd2 * ((2'd2)&&(2'd3))));
  localparam [5:0] p14 = ((2'd1)?(3'sd3):(&(5'd8)));
  localparam signed [3:0] p15 = (5'sd11);
  localparam signed [4:0] p16 = {(4'd14),(2'd0),(2'd1)};
  localparam signed [5:0] p17 = ({1{(((4'sd6)?(3'd7):(5'sd7))!==((-5'sd5)&(5'd7)))}}?{{2{(4'd0)}},{3{(-4'sd3)}},{2{(5'd0)}}}:{1{{1{{3{(3'sd1)}}}}}});

  assign y0 = {(5'd17),$signed((a4?a0:a3))};
  assign y1 = {((~|(p15?p13:b2))^{(p0?p16:p11)}),{(~^(4'd2))}};
  assign y2 = ((b5?b1:a5)?(a3?b0:p14):(b3?b0:a4));
  assign y3 = $signed((((p16?a0:b4)<<<(+b0))?((~^a2)%p5):$signed((a5<<a3))));
  assign y4 = ($unsigned((b2<p8)));
  assign y5 = (-5'sd2);
  assign y6 = (!(&(((~^(^(-5'sd0)))!=((|a3)>>(^b5)))^((+(-4'sd6))|(-2'sd1)))));
  assign y7 = (((b0?p11:b0)<=(3'sd1))?({b1,a3}>=(b5!==a0)):((3'sd0)?(~&a3):(4'd2 * b1)));
  assign y8 = $signed($unsigned($unsigned($unsigned((&((-((p9^a2)&(b1)))<={3{{2{p5}}}}))))));
  assign y9 = (~^((-2'sd1)<<<(3'd4)));
  assign y10 = ({(&a0)}?(&(-b3)):(p7==p6));
  assign y11 = (~|{2{(b1?b1:a3)}});
  assign y12 = {(((p12==a3)&(|(-b2)))!=({b0,a5,p3}!={(5'sd4)}))};
  assign y13 = ({(b1<b5)}?(a2!=p6):{(a5&p1)});
  assign y14 = (a2>>a1);
  assign y15 = (2'sd0);
  assign y16 = $unsigned({(b5+a2),(b2===a3),$signed(b0)});
  assign y17 = {1{((~(5'd2 * b1))=={2{(~^b4)}})}};
endmodule
