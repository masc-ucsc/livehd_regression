module expression_00701(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(-5'sd2),(4'sd5),(-4'sd5)},(&((-4'sd2)?(2'd1):(4'sd2))),((2'd1)?(2'd0):(3'd6))};
  localparam [4:0] p1 = {1{{{1{{3{(2'sd0)}}}},{((4'd15)?(5'd19):(5'd16))},((2'd3)<<<(3'd2))}}};
  localparam [5:0] p2 = ((-5'sd14)<=({3{(3'sd2)}}<<<((-2'sd0)!=(-4'sd5))));
  localparam signed [3:0] p3 = ({4{(~&(2'd1))}}>((6'd2 * (4'd12))?((-5'sd6)?(4'd15):(3'd2)):(|((-2'sd0)<<<(4'sd2)))));
  localparam signed [4:0] p4 = (2'sd0);
  localparam signed [5:0] p5 = {2{(((5'd31)?(-4'sd3):(4'sd4))?((5'sd0)?(4'sd0):(-4'sd1)):(4'd2 * (5'd31)))}};
  localparam [3:0] p6 = (((4'd7)<=(4'd1))?((4'd3)?(2'd1):(5'sd3)):((5'd25)||(2'd2)));
  localparam [4:0] p7 = (((&{(4'd3)})-((4'sd4)+(4'd4)))>=(~{(~^(5'sd13)),{(3'sd1)},(!(4'sd3))}));
  localparam [5:0] p8 = (!(2'd0));
  localparam signed [3:0] p9 = (5'd0);
  localparam signed [4:0] p10 = {(~|(3'sd0)),{1{(4'sd0)}}};
  localparam signed [5:0] p11 = (((3'd4)?(3'd3):(4'd10))?(+(2'd0)):{4{(2'sd1)}});
  localparam [3:0] p12 = (((5'd2)<=(2'd1))?(5'd18):((4'd2)===(3'd0)));
  localparam [4:0] p13 = {3{(4'd9)}};
  localparam [5:0] p14 = (-4'sd3);
  localparam signed [3:0] p15 = ((+(((-3'sd2)|(3'd7))%(4'd2)))>((|((2'd2)*(3'd2)))<<(&((4'd11)==(-3'sd0)))));
  localparam signed [4:0] p16 = {3{(!{4{(2'sd1)}})}};
  localparam signed [5:0] p17 = {2{((5'd2 * (5'd29))<((3'd6)>=(5'd21)))}};

  assign y0 = {3{((p17&p1)!=(^b0))}};
  assign y1 = $unsigned(a5);
  assign y2 = ((5'sd6)?(~|p8):(p0?p2:p0));
  assign y3 = {(-2'sd1),{{a5,p4,b4}},(~&(-2'sd0))};
  assign y4 = (~^(|((~^(a1&&a5))>>((~|b2)+(a2?a5:p13)))));
  assign y5 = {3{{1{p16}}}};
  assign y6 = ($unsigned({{({a5,p1,p11}?(a0?a5:p7):{2{p12}})}})|((((5'd9)>>>(b3>b2)))!=={4{b4}}));
  assign y7 = ((p17>>p11));
  assign y8 = {({b1}?{2{a5}}:{b4,p3,p7}),(+$signed($signed({2{p2}})))};
  assign y9 = ((b5>=b4)<(-2'sd0));
  assign y10 = (-5'sd7);
  assign y11 = ((p16%b5)%b4);
  assign y12 = ((-(|$signed(b4)))^(+$unsigned($signed(p15))));
  assign y13 = $signed($signed((p16?a4:a3)));
  assign y14 = ((-(2'd0))<=((b2&&b2)>>>$signed((2'd0))));
  assign y15 = {2{(~&({a5}>{p6,p13,p10}))}};
  assign y16 = (^(^(~|{2{(!$unsigned($unsigned(((b3<<a1)<<<(a3+p5)))))}})));
  assign y17 = (4'd13);
endmodule
