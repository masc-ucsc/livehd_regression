module expression_00075(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd9)^(5'd13))^~((-3'sd0)?(5'sd12):(3'd2)));
  localparam [4:0] p1 = {(2'd0),(-2'sd1),(5'sd14)};
  localparam [5:0] p2 = ((|(((2'sd1)!==(4'd14))===((5'sd3)*(2'sd1))))?(((-3'sd0)||(-4'sd0))?((3'd4)%(4'd3)):(^(2'd3))):((~|(-3'sd0))<=((5'd6)?(5'd30):(-3'sd0))));
  localparam signed [3:0] p3 = (!({((~|(3'd3))!=((-2'sd0)&&(4'd9)))}>=(5'd2 * (~&{(3'd5)}))));
  localparam signed [4:0] p4 = (~^(&(~&(~&(~^(~((4'd4)^~(4'd3))))))));
  localparam signed [5:0] p5 = {{(2'sd1)}};
  localparam [3:0] p6 = ((+(2'd0))?(((2'd3)?(2'sd0):(4'sd1))^((2'sd0)?(-5'sd12):(2'sd0))):((3'd3)?(3'd1):(-3'sd1)));
  localparam [4:0] p7 = (({1{(5'sd1)}}?{(-2'sd1),(2'sd0),(5'd1)}:((-3'sd2)|(-4'sd2)))?(((3'd1)?(-4'sd3):(-3'sd1))^((3'd4)&(2'd1))):({2{(-4'sd6)}}?((2'd2)==(5'sd12)):{(-3'sd0),(2'd2)}));
  localparam [5:0] p8 = {2{(|{1{(2'sd0)}})}};
  localparam signed [3:0] p9 = (-{4{(3'd6)}});
  localparam signed [4:0] p10 = ({(-3'sd0),(3'd4)}|((2'd0)?(2'd2):(3'd2)));
  localparam signed [5:0] p11 = (3'd6);
  localparam [3:0] p12 = (((&((-5'sd7)>>(-5'sd1)))&((5'sd13)?(5'sd13):(-2'sd0)))>>(~&(&(+((~^(2'd3))-(|(3'd5)))))));
  localparam [4:0] p13 = ((5'd10)===(3'd0));
  localparam [5:0] p14 = (((4'sd0)|(3'd4))-((2'd2)!=(5'd22)));
  localparam signed [3:0] p15 = (4'd6);
  localparam signed [4:0] p16 = {(-3'sd0),(-4'sd0),(5'd2)};
  localparam signed [5:0] p17 = ({(&(-(3'd2))),{2{(4'd10)}},{3{(2'sd1)}}}=={{1{(+{{(2'd3)},((-2'sd1)||(2'd0))})}}});

  assign y0 = (4'd2 * (p14+a1));
  assign y1 = (-({4{(a5-b3)}}?((~|(p1))^(b0?p14:p1)):((4'sd3)>=$unsigned($unsigned(b1)))));
  assign y2 = ((((~|(~|p13))&(3'sd0)))^~$signed({{p1,p15,p12},(p8^~p6),(|a5)}));
  assign y3 = ((|(+(p9&b2)))>>(2'd3));
  assign y4 = {{(({p5,p5,p3}^((a5)===(5'd23))))}};
  assign y5 = {3{$unsigned(({2{p10}}))}};
  assign y6 = (5'd2 * $unsigned($signed(p15)));
  assign y7 = (-$unsigned((($signed((-{b3,p3,a2}))+(!(b2===a3)))&&(2'd0))));
  assign y8 = (+{(~({p4,a1}>>>{p16,p4,a1}))});
  assign y9 = ((-{(b4),(-p1),(p0<<a5)})>$signed($unsigned((~^$signed({(b2)})))));
  assign y10 = {(p13<=p3),$signed({p8,b3}),(a5!=a2)};
  assign y11 = (p3||p3);
  assign y12 = ({(^$unsigned(($unsigned((((b0>>p9)<<(~^{p7,p10}))<<<(((p4!=p16)|((a5===a5)))))))))});
  assign y13 = $signed((~|(^(~^p13))));
  assign y14 = (2'd1);
  assign y15 = (((p2?b5:b3)?(a3?p2:p11):(&p0))?(^(-((~b3)?(+a1):(~^p6)))):(|(~((p2?p10:a3)?(p8?p14:p0):(a1?p1:b3)))));
  assign y16 = (((^(+(~p13)))!=((a5&&p0)<=(p14^a4)))!=(4'd2 * (p14<=p13)));
  assign y17 = ((p6%p14)||(b3|p13));
endmodule
