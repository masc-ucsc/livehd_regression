module expression_00057(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'sd2)?(3'sd2):(4'd12));
  localparam [4:0] p1 = (5'd2 * ((5'd25)<<(3'd5)));
  localparam [5:0] p2 = ({3{(2'sd0)}}<<((3'd7)>(3'd6)));
  localparam signed [3:0] p3 = {{3{(5'd16)}},{((-5'sd15)?(4'sd0):(2'd0))},((2'sd0)!=(5'd4))};
  localparam signed [4:0] p4 = ((2'd3)||(-4'sd1));
  localparam signed [5:0] p5 = (5'sd3);
  localparam [3:0] p6 = {4{(-2'sd1)}};
  localparam [4:0] p7 = ((((2'd0)?(4'sd2):(4'sd1))==(5'sd5))===(4'sd6));
  localparam [5:0] p8 = (!(!{2{((4'd0)?(5'd0):(3'sd0))}}));
  localparam signed [3:0] p9 = {3{(((2'sd0)^~(5'd20))>((-3'sd0)>>(4'sd2)))}};
  localparam signed [4:0] p10 = (-(+{3{(~&(~&(5'sd5)))}}));
  localparam signed [5:0] p11 = {3{(((-5'sd14)&(3'd2))?((2'd2)>(-5'sd2)):((2'd3)!==(4'sd3)))}};
  localparam [3:0] p12 = (5'sd1);
  localparam [4:0] p13 = ({(5'd26),(-4'sd3),(2'sd0)}&&((4'sd5)==(2'sd0)));
  localparam [5:0] p14 = ({((-3'sd2)!==(-3'sd2)),{4{(3'd7)}},{(4'd13)}}?({3{(2'd1)}}?((2'd3)>(3'd5)):((3'd5)!=(-3'sd2))):((5'd6)>=(!(4'd10))));
  localparam signed [3:0] p15 = ((-2'sd0)|(2'sd1));
  localparam signed [4:0] p16 = (~^(~(~^(3'd6))));
  localparam signed [5:0] p17 = (((~|(-3'sd3))&((4'd1)?(5'd11):(5'd18)))?((4'sd2)?(3'd4):(4'sd0)):(((-3'sd1)&&(4'd11))<<{1{(2'd0)}}));

  assign y0 = (((b4|a0)-(6'd2 * b1))&((a2===b2)|(a2>>>p10)));
  assign y1 = ((~&$unsigned($unsigned($signed((-((~{1{$signed($unsigned({3{$signed(b1)}}))}}))))))));
  assign y2 = (!(a0!=a5));
  assign y3 = {1{{3{(2'd1)}}}};
  assign y4 = ((-3'sd3)-(2'd0));
  assign y5 = ({$signed(a2),(&b2)});
  assign y6 = (-2'sd1);
  assign y7 = ($unsigned(((~b1)))?(~^$signed({b3,p10,p17})):{p0,a1,b0});
  assign y8 = (-(!($signed({3{p9}})<(p4?b4:b5))));
  assign y9 = ((6'd2 * a1)?(b3?p15:a1):(p10?p2:b0));
  assign y10 = (((b2===b5)?(p8^~p2):(b3!=b4))?((p1?p13:p15)?(b5*b1):(b4!=b5)):((b2>a4)^(a1<p14)));
  assign y11 = ((((b3&&a2)>>(b5))));
  assign y12 = {(-2'sd0),(3'sd2)};
  assign y13 = ({(b4>>>a4)}?(+(-2'sd1)):(^(a0===b4)));
  assign y14 = $unsigned(((!(b1?a0:a2))?{2{(a0)}}:(-3'sd1)));
  assign y15 = (4'd6);
  assign y16 = $unsigned((~|{3{($unsigned(p9)!=$signed(a0))}}));
  assign y17 = (((b2<<a4)+{a4})===((!a0)||(a4+a3)));
endmodule
