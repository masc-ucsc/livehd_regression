module expression_00869(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{{(5'd15),(5'd5),(3'd5)}}};
  localparam [4:0] p1 = ({4{(3'd5)}}>((2'd1)>(-4'sd3)));
  localparam [5:0] p2 = {{(2'd1),(2'd2),(4'sd4)},(+{(5'sd9),(5'd30),(-5'sd5)}),{{(3'sd2),(3'd5)}}};
  localparam signed [3:0] p3 = {1{{({4{(2'd1)}}|((-5'sd7)>=(3'sd1))),(~{{1{(5'sd7)}},{3{(-2'sd1)}}})}}};
  localparam signed [4:0] p4 = (5'd2 * {(~(3'd6))});
  localparam signed [5:0] p5 = (!((((5'd2)!==(-5'sd12))&&(3'd2))&(&(2'd3))));
  localparam [3:0] p6 = ((~&((4'd7)?(3'sd1):(3'sd0)))?{{(-3'sd3),(2'sd1),(-4'sd4)}}:(~&(3'd6)));
  localparam [4:0] p7 = (~&((&(&(-(2'sd0))))?(|(+((5'd19)?(5'd20):(3'd3)))):(-{1{(5'd6)}})));
  localparam [5:0] p8 = {{3{(5'sd10)}},{4{(2'd1)}}};
  localparam signed [3:0] p9 = (|(&{(&((((5'd20)?(-2'sd0):(5'sd11))||((2'sd1)>(3'd0)))!==(((2'd2)!=(5'sd13))?(~|(5'd11)):{(3'd4)})))}));
  localparam signed [4:0] p10 = (~&(-5'sd8));
  localparam signed [5:0] p11 = (5'd18);
  localparam [3:0] p12 = ((((-5'sd7)^~(2'd3))!==((2'd1)<=(5'd30)))&((2'sd1)^((4'd14)?(5'sd12):(4'd5))));
  localparam [4:0] p13 = ((-3'sd3)?(&(&(2'd2))):(^(&(-2'sd0))));
  localparam [5:0] p14 = (~^(-5'sd6));
  localparam signed [3:0] p15 = (5'd10);
  localparam signed [4:0] p16 = ((((3'sd0)?(2'd2):(3'sd2))?((3'sd3)<(3'd6)):((4'sd3)||(-2'sd0)))>>(((5'd7)?(-3'sd0):(2'd2))&&((-5'sd12)&(-4'sd7))));
  localparam signed [5:0] p17 = ({4{(4'sd6)}}!=(~^(!(-2'sd0))));

  assign y0 = (2'sd1);
  assign y1 = (a3!==a2);
  assign y2 = (~b5);
  assign y3 = $unsigned(((((a5)?(p10?p6:p7):(a0<a3))<$signed((p16?b2:p11)))));
  assign y4 = (+(!((+(&(({2{b1}}||(b5?b5:a4))?({2{b5}}?(b1<<<b1):(-a2)):({3{a1}}!=(+b1))))))));
  assign y5 = ((-(&((^(b4<<b3))^~(a1?a3:b0))))===({2{b2}}?(a4?a2:b2):(a4?b3:a2)));
  assign y6 = (&((a3>=a0)*(a1>>a5)));
  assign y7 = ($unsigned((3'd3))?(2'd1):(~&((p9<<a5)!=(p9?p4:a1))));
  assign y8 = {1{{1{(b4-b2)}}}};
  assign y9 = {1{(~((!{4{(b0^b4)}})!=={3{{4{a5}}}}))}};
  assign y10 = ((p14?b2:p9)?(p13+p11):(p17?p17:p8));
  assign y11 = {{3{{1{b5}}}},{{1{p12}},{1{p0}}},{(a0),{a4,b2}}};
  assign y12 = {{{(!(b2<<<b1))},({1{b0}}>>>(2'd1))},(~&(~^((4'sd7)|(&(b0|a4)))))};
  assign y13 = (({b2,p0,p0}?(p9?a0:p3):(+p2))?{(~p2),{p10,p14}}:(~(~{(~^a1)})));
  assign y14 = {((5'd5)?{(p12?p0:p9),(a2===a1)}:({4{b1}}==(p13||p6)))};
  assign y15 = (^(((a4===b5)!==(+(b1>a3)))>>>({1{{3{p13}}}}|(p4<=p2))));
  assign y16 = (|(~$unsigned((&(~&(~^{2{((6'd2 * p6)!={b2,b4,a3})}}))))));
  assign y17 = $signed((((a1!=b0)?{1{a0}}:(a3<a3))?({1{(6'd2 * a2)}}-(-(3'sd2))):(-4'sd4)));
endmodule
