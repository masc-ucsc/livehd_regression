module expression_00714(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd30);
  localparam [4:0] p1 = {{{(4'd13),(3'd7)},((2'd1)?(4'd0):(3'd4)),(!(5'd30))},{2{((5'd16)||(3'd1))}}};
  localparam [5:0] p2 = (~&(5'd22));
  localparam signed [3:0] p3 = {2{(-(((2'd3)&(4'd15))?(~&(4'd4)):{2{(2'sd0)}}))}};
  localparam signed [4:0] p4 = ((5'd19)||(-4'sd7));
  localparam signed [5:0] p5 = ({3{((2'sd1)!=(2'd0))}}==(|(~&(~((5'sd5)<<<(4'sd3))))));
  localparam [3:0] p6 = (5'd6);
  localparam [4:0] p7 = {(&{(5'd2)}),{3{(3'd1)}},((-4'sd2)!=(5'd5))};
  localparam [5:0] p8 = (3'sd1);
  localparam signed [3:0] p9 = (-(~^(~(~^(2'd1)))));
  localparam signed [4:0] p10 = (2'd2);
  localparam signed [5:0] p11 = (5'd11);
  localparam [3:0] p12 = ({(4'sd5),(5'd17)}?(5'd5):{(-5'sd14),(5'sd4)});
  localparam [4:0] p13 = ((((2'sd1)>>>(5'd11))^((-5'sd4)?(5'd7):(-2'sd1)))!==((3'd7)>=((-3'sd2)>(2'd2))));
  localparam [5:0] p14 = ((|(4'd2 * ((3'd4)/(5'd19))))>((-4'sd3)^~(2'd1)));
  localparam signed [3:0] p15 = {(2'd1),(-2'sd0)};
  localparam signed [4:0] p16 = ((((-3'sd1)>(4'sd4))^~((4'd11)&(2'd2)))^~(((-3'sd0)<<<(-5'sd1))+((3'sd0)^(5'd6))));
  localparam signed [5:0] p17 = (~^{(3'sd2),(5'd27)});

  assign y0 = (4'd5);
  assign y1 = {(~|(p11-b1)),{1{{p17,a5,b0}}},(~^(5'sd7))};
  assign y2 = {(&{4{p2}}),(~(b1|p5)),$unsigned($unsigned(p13))};
  assign y3 = (|a4);
  assign y4 = ({3{b1}}?{4{a4}}:(p5?p1:a3));
  assign y5 = {2{{2{(-(~^p6))}}}};
  assign y6 = {(~&{{(!b0),{b2,a1}},(+(!{b1,a5})),{p11,a1,a5}})};
  assign y7 = (p15?p16:p4);
  assign y8 = (((&b4)?(~|a3):(a5?a2:b5))?(~^(b5?p16:a2)):((b5<<b5)|(a1<p17)));
  assign y9 = (((-4'sd6)%a1)>((3'd0)+(3'd2)));
  assign y10 = (((5'd2 * p12)^~(6'd2 * p6))?((a0|p7)^(p17|p17)):((p3^~p17)?(p14^p0):{a3,p12,p15}));
  assign y11 = ((a5||a2)+{4{b1}});
  assign y12 = {{b3,b5,p1},{a5,a0,a3},(-5'sd1)};
  assign y13 = (((p13?b0:p0)?(5'sd5):(b4>p5))?((b5?p5:p12)?(a5?p1:p2):(a4+a5)):((p11?p4:p11)?(p16>p13):(p17/p3)));
  assign y14 = (b1^~p0);
  assign y15 = (3'd6);
  assign y16 = {p13,p16,b0};
  assign y17 = (((!b1)?(a4?p8:a3):(~b3))?(+(~|(~(~^(~^a0))))):(-2'sd0));
endmodule
