module expression_00720(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'd11);
  localparam [4:0] p1 = ((((-3'sd0)?(2'd0):(-3'sd2))>{(2'd3),(2'd1)})>>(((3'd5)<=(5'd14))!={(2'sd0),(3'd3)}));
  localparam [5:0] p2 = (+(&(4'd4)));
  localparam signed [3:0] p3 = ((^(~^(5'sd10)))&(~|(&(4'd3))));
  localparam signed [4:0] p4 = {3{{3{(5'd3)}}}};
  localparam signed [5:0] p5 = {3{(3'sd2)}};
  localparam [3:0] p6 = ({{(~^(-5'sd3))},(^{(5'sd2),(2'd3)})}>{((3'sd0)===(5'd1)),{(2'd3)},(~^(3'd3))});
  localparam [4:0] p7 = (-(|(-(|(-((4'd0)>>>(3'sd2)))))));
  localparam [5:0] p8 = ({(-5'sd3),(5'd4)}?{(5'd17),(-3'sd1)}:((-4'sd0)==(2'sd0)));
  localparam signed [3:0] p9 = {(5'd10),(5'sd14)};
  localparam signed [4:0] p10 = ({{{(-2'sd1)}},((4'd9)^~(3'd4)),((2'sd0)<<<(3'd5))}&&(((2'd3)||(4'd2 * (5'd2)))!=(2'd0)));
  localparam signed [5:0] p11 = (|({(3'd3),(-3'sd1)}<<<(-4'sd6)));
  localparam [3:0] p12 = ((^(2'd1))!==(5'd2 * ((2'd2)>=(2'd3))));
  localparam [4:0] p13 = ((~((+(4'd1))<<(~^(-2'sd0))))>>>(&(-(&((~|(-2'sd0))<<<((2'd2)<<(-3'sd2)))))));
  localparam [5:0] p14 = (5'd15);
  localparam signed [3:0] p15 = (^(!((((5'd0)>>>(-5'sd12))<=(&(5'd2 * (3'd4))))&(|{1{{{2{(4'd11)}},{(3'd4),(4'd11),(2'sd0)},((2'sd0)>(-3'sd3))}}}))));
  localparam signed [4:0] p16 = ((4'd12)<<<(5'd7));
  localparam signed [5:0] p17 = (4'sd2);

  assign y0 = ((+(~|(^(+(~|(^(~^(p13>>p14))))))))>=(|(^((~^(~&p6))||{2{a2}}))));
  assign y1 = ((-((~(b1>>>a1))-(b0<=a5)))||(~|((~|(p12&&b0))%a5)));
  assign y2 = (!(-b3));
  assign y3 = {2{(+(|(-$unsigned(((+((-(~|b4)))))))))}};
  assign y4 = (((a5==p1)?(a0>=p11):(b0<<p13))||(~^((a5?p5:p16)>>>(b5<<<a0))));
  assign y5 = ((($unsigned(p4)?(p8||p9):{3{p17}})<(+((|(p9==p14))>>>$unsigned((p14^p11))))));
  assign y6 = {{({a2,a2,b5}!==(~{a1}))}};
  assign y7 = $unsigned(((~|{4{p0}})+((3'sd3)?(p2&p17):(p6>p4))));
  assign y8 = (((b0<=a1)^~(a5<=a4))|((a1%a1)&&(a4!=a0)));
  assign y9 = (~^$unsigned(({(a2+a3),{b2,b4},{b3,a1,b1}}<<<(&(~^{b5,a2,b1})))));
  assign y10 = ($unsigned({(+a0),(b0?a1:a0)})?(~^{{(a1)}}):$unsigned((a4?a3:b3)));
  assign y11 = {(4'd8),{(~(4'd0))}};
  assign y12 = $unsigned(($signed(p5)?(b3):(a5?b3:b4)));
  assign y13 = {4{{4{a0}}}};
  assign y14 = ((&{4{p13}})&&({p13,p9,p13}>>(^a5)));
  assign y15 = (((5'd2 * a0)<=(p0!=b4))?((b1)!=(~&p2)):((p12?p11:p11)));
  assign y16 = (~&(&(~^(^(^(~&((|(-2'sd1))?(2'd2):(a4?b5:a5))))))));
  assign y17 = (5'd3);
endmodule
