module expression_00993(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((2'd0)?(2'sd0):(5'sd8)),{(-2'sd1),(-2'sd0)},(+(-2'sd1))};
  localparam [4:0] p1 = ((4'd13)<=(-2'sd1));
  localparam [5:0] p2 = (({2{((-4'sd0)!==(3'sd3))}}-(((3'sd2)<<(-3'sd1))==(2'd3)))>>({1{(~|((2'sd1)==(4'd5)))}}!=(((4'd10)===(-2'sd1))<<<((3'sd3)>>>(3'sd2)))));
  localparam signed [3:0] p3 = ((2'd2)<<(3'd1));
  localparam signed [4:0] p4 = (5'd4);
  localparam signed [5:0] p5 = ((-{4{(3'sd3)}})<<((3'sd0)+(-5'sd13)));
  localparam [3:0] p6 = ({2{((2'd1)!=(5'sd1))}}!=(^({3{(3'd3)}}!={(4'sd6),(4'd2),(2'd2)})));
  localparam [4:0] p7 = (|(~&(~^(&(~&(~(5'sd12)))))));
  localparam [5:0] p8 = ({(|((3'd4)^~(3'd5)))}-((2'd3)?(3'sd3):(4'd11)));
  localparam signed [3:0] p9 = (3'sd1);
  localparam signed [4:0] p10 = (2'd1);
  localparam signed [5:0] p11 = (4'sd2);
  localparam [3:0] p12 = ((4'd11)==(3'sd2));
  localparam [4:0] p13 = (4'd9);
  localparam [5:0] p14 = (((-3'sd0)?(3'sd2):(3'd7))?((3'sd1)?(3'd1):(4'sd5)):(+(4'd8)));
  localparam signed [3:0] p15 = ((2'd1)?({4{(4'd9)}}?((4'd2)?(2'sd1):(5'd13)):{(-4'sd5),(5'd10),(2'd1)}):{((2'd0)?(5'd15):(2'sd0)),((-5'sd11)<(3'd5))});
  localparam signed [4:0] p16 = (((5'd30)==(3'd7))<=((-3'sd2)!==(4'sd1)));
  localparam signed [5:0] p17 = ((3'd5)?(3'd2):(3'd6));

  assign y0 = (~&{{p11,a0,p1},(p6?p4:a4)});
  assign y1 = (&((-p2)<<(p14)));
  assign y2 = {1{{1{(((a4&&a3)===(a5&&b5))>>{3{(a2==a5)}})}}}};
  assign y3 = ({((~^p7)?(p8?p4:p4):(~|p14)),(((p5<<p10)<<<$unsigned(p14))),((p12||a0)^~(p7<<<p0))});
  assign y4 = (((p2?b4:b4)?(p11?p0:b3):(b2?a5:a4))?((p10?p2:p1)?(b4?a3:b0):(a4?a5:b0)):((b1?p9:b1)?(p1?b4:a2):(a2?p2:p7)));
  assign y5 = (^{(5'd2 * p6),(~^a3),{3{p0}}});
  assign y6 = $unsigned($unsigned($unsigned((^(~((a1!==a3)%p4))))));
  assign y7 = ($signed({({2{p1}}?{4{p3}}:{1{p11}})})&{(&{p7,a1}),{$signed({1{p11}})}});
  assign y8 = {2{{4{(a5>=b2)}}}};
  assign y9 = (-5'sd13);
  assign y10 = {(5'd2 * (a1>=p6))};
  assign y11 = (a0?p5:p9);
  assign y12 = (+(^(&a4)));
  assign y13 = (~^((-4'sd7)^(p13^p12)));
  assign y14 = (((b5^~b3)<=$unsigned(a5))^{(a3<<<a2)});
  assign y15 = {1{{2{($signed((b0-a1))|($unsigned(a3)^~(p8?b1:a2)))}}}};
  assign y16 = (p10|p13);
  assign y17 = $signed((((p16?a5:b5)?(2'd1):$unsigned((b0)))&&$signed((6'd2 * {4{a2}}))));
endmodule
