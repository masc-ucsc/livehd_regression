module expression_00201(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd15);
  localparam [4:0] p1 = ((((2'd2)<(-3'sd3))?((-4'sd3)>>(5'd28)):(!(5'sd13)))?(((5'd24)<(5'd6))?((-4'sd1)!==(4'd14)):(6'd2 * (2'd1))):(((-5'sd6)+(-3'sd0))+((2'd0)>>(4'sd1))));
  localparam [5:0] p2 = ((3'd3)*(5'd10));
  localparam signed [3:0] p3 = (~&((!((4'd1)<<(3'd4)))<<(^((5'd4)|(5'd26)))));
  localparam signed [4:0] p4 = (^(!((^(+(|((5'd30)&(4'd3)))))&((!(3'sd0))>(^(5'd9))))));
  localparam signed [5:0] p5 = {({(-3'sd3)}||{1{(4'd7)}}),(((5'd20)^~(-5'sd1))||(!(-5'sd1)))};
  localparam [3:0] p6 = (!(+(2'd0)));
  localparam [4:0] p7 = ((5'd30)<((-4'sd5)|(2'd3)));
  localparam [5:0] p8 = (+(5'd31));
  localparam signed [3:0] p9 = {1{{2{(-3'sd0)}}}};
  localparam signed [4:0] p10 = {2{((-5'sd8)?(4'sd7):(3'd3))}};
  localparam signed [5:0] p11 = {1{((((2'd0)|(5'd6))!==((5'sd12)&(3'sd2)))=={4{(5'd27)}})}};
  localparam [3:0] p12 = (|((-3'sd2)>>>(2'd3)));
  localparam [4:0] p13 = {1{(!(((2'sd0)<<(3'd7))<<(-{4{(2'd0)}})))}};
  localparam [5:0] p14 = (((3'sd2)-(-2'sd1))+{4{(5'd12)}});
  localparam signed [3:0] p15 = (((6'd2 * (5'd7))!==((4'd4)!==(5'sd15)))^(((-5'sd5)==(3'd0))=={(3'sd0)}));
  localparam signed [4:0] p16 = (-5'sd7);
  localparam signed [5:0] p17 = (!(4'd12));

  assign y0 = ((a0===a1)>(p0&&p17));
  assign y1 = {1{(-3'sd0)}};
  assign y2 = (+((a4?b0:a4)!==$unsigned((a3?a3:b2))));
  assign y3 = (({2{a3}}!=(b3?b1:b5))-((a4===a5)<(a1^a0)));
  assign y4 = (~(b3===b0));
  assign y5 = ((((!(|a2))%b0)^(~|((~^a2)%a0)))<((|(~&(a2==a1)))==((6'd2 * b1)&(~|a1))));
  assign y6 = (a4^b2);
  assign y7 = ((^((~|{p5,b5})))>>$unsigned((~&(b1?p6:p13))));
  assign y8 = {(((a4||p12)?(~^(p16^p1)):(|(a2===b5))))};
  assign y9 = ((2'd2)?(b0?p9:p1):(p3?p0:p14));
  assign y10 = {2{{{2{p9}}}}};
  assign y11 = ((|(!(+(p12&&p3))))<=(~^((p1==p8)*(|b2))));
  assign y12 = (((p14?a1:b1)?(&p14):{4{p16}})?((p14>p7)<<{b1,b5,b5}):(^{{4{p1}},(+b2)}));
  assign y13 = (a2<=p14);
  assign y14 = ((~((+(!b1))>>{3{b4}}))!=={4{{a5,b1}}});
  assign y15 = (((~&p1)!=(p7>>>p7))?({p11,p12,p3}<<<(p8?p11:p11)):(p16?p0:p17));
  assign y16 = $unsigned((|{4{(4'sd5)}}));
  assign y17 = (~&$unsigned((({4{a1}}!=={2{$signed(a0)}})>>>{2{$unsigned((p7-p11))}})));
endmodule
