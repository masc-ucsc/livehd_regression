module expression_00023(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{((2'd1)?(2'd1):(2'd2))}};
  localparam [4:0] p1 = {((5'd10)!=(~|{(3'sd1),(3'd1),(4'd3)}))};
  localparam [5:0] p2 = ((2'd0)|(2'sd1));
  localparam signed [3:0] p3 = (-4'sd1);
  localparam signed [4:0] p4 = {1{(~^((~|(5'sd9))?((-3'sd0)?(5'd10):(5'd28)):(|(2'd2))))}};
  localparam signed [5:0] p5 = {3{{2{(3'sd0)}}}};
  localparam [3:0] p6 = (4'd8);
  localparam [4:0] p7 = (|(^{(-3'sd1),(-2'sd0),(2'd2)}));
  localparam [5:0] p8 = {2{({2{((4'd9)?(3'd0):(4'd10))}}^~{1{{3{(5'sd7)}}}})}};
  localparam signed [3:0] p9 = (|(-(((5'd18)>=(5'sd9))*((5'd9)<<(3'd6)))));
  localparam signed [4:0] p10 = (&((4'd12)/(5'd25)));
  localparam signed [5:0] p11 = (+{(-{1{(-3'sd2)}}),{(~^(3'd0)),(~^(6'd2 * (5'd9)))}});
  localparam [3:0] p12 = ((((-3'sd2)&&(3'sd1))<{(4'd8),(3'd6)})<=(((3'd4)^(4'sd7))+((-4'sd1)|(2'sd0))));
  localparam [4:0] p13 = ((~|((5'd24)?(-5'sd10):(-3'sd1)))?(-5'sd3):(!(~^((3'd6)>(4'd12)))));
  localparam [5:0] p14 = (-2'sd1);
  localparam signed [3:0] p15 = (((5'd4)===(-5'sd12))>>>{3{(-2'sd1)}});
  localparam signed [4:0] p16 = (-(-(4'sd5)));
  localparam signed [5:0] p17 = (5'd2 * (&(~(5'd31))));

  assign y0 = {{(a1===b1),{1{(^a4)}}},{2{(4'd2 * b1)}},((-(~&a0))!=={2{a1}})};
  assign y1 = {(^$signed({{(a5),(~^a0),$signed(a0)},({a5,b4,a0}>(b3>=a2)),{((b1)!=(+b3))}}))};
  assign y2 = ({($signed(((b1<<p16)<=(3'd3)))^(2'd1))});
  assign y3 = ({1{(-((6'd2 * p1)^(|(^p16))))}}-(!((~|p13)?(p15>>>p0):(!p9))));
  assign y4 = {p15};
  assign y5 = (~((&p4)<<(|p14)));
  assign y6 = (({4{a0}}+({3{a4}}<<(3'd1)))>{4{{3{a1}}}});
  assign y7 = ({4{{2{{2{p10}}}}}});
  assign y8 = (-2'sd1);
  assign y9 = ({((b3+a4)?{a1,b1,b5}:(b5>=p14))}|{(b0<<a0),{(b3?a5:p13)}});
  assign y10 = $unsigned((((a0==a4))?(^(b5)):(a0?a2:p3)));
  assign y11 = {4{(^{1{(+(~|p7))}})}};
  assign y12 = ((b2>>a4)?(a5?p9:b5):{1{p11}});
  assign y13 = {3{{3{p17}}}};
  assign y14 = (|{(~|({p1,p0,p6}|(+p0))),(~&{(p1>>p17)}),((~p6)<=(+p5))});
  assign y15 = (^(~|(!{2{(~p8)}})));
  assign y16 = {{(~((p9&&p4)==(^(a5>b5))))}};
  assign y17 = (~^(~&(p9<=p4)));
endmodule
