module expression_00713(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd1);
  localparam [4:0] p1 = {(+{((~^(-5'sd0))?(&(5'd25)):{(-3'sd1),(3'd0)}),{((2'd3)?(3'd1):(4'd10)),((3'd7)?(5'd17):(3'd3)),(5'sd5)}})};
  localparam [5:0] p2 = (~^((((3'd5)&&(5'd20))||{(2'sd1),(3'd0)})==(4'd3)));
  localparam signed [3:0] p3 = (~^(~&(~|(+{1{(~&(((-3'sd2)-(4'd15))==(|(&(5'sd1)))))}}))));
  localparam signed [4:0] p4 = (~|{(((2'd2)>>>(3'sd0))>=(|(2'sd1))),(&(5'd2 * (4'd5)))});
  localparam signed [5:0] p5 = ({{4{(-2'sd1)}}}?(|((4'd12)|(-4'sd3))):((5'd3)&&(5'd3)));
  localparam [3:0] p6 = (2'd1);
  localparam [4:0] p7 = ({3{(4'd13)}}>>>((3'd4)<=(3'sd0)));
  localparam [5:0] p8 = (((~(5'd2 * (2'd2)))==={((-4'sd3)^(2'd3))})&{((4'd11)<<(-2'sd0)),((4'd15)&&(-2'sd0))});
  localparam signed [3:0] p9 = (((3'sd3)+(2'sd1))<((4'd7)>>>(2'd0)));
  localparam signed [4:0] p10 = ((((-2'sd0)?(5'd25):(-4'sd6))?(4'sd2):((4'sd5)?(2'd2):(-5'sd5)))?(-5'sd6):(((2'd0)?(2'sd1):(3'sd3))?(5'd27):(-5'sd14)));
  localparam signed [5:0] p11 = (!(~({(2'd2),(2'd3),(4'sd4)}==(-2'sd1))));
  localparam [3:0] p12 = (2'sd0);
  localparam [4:0] p13 = {{{3{(2'sd1)}},{1{{(3'sd3),(2'sd1),(5'd14)}}}},(|({(2'd1),(2'd0),(3'd4)}>(4'd6)))};
  localparam [5:0] p14 = ({(4'd0),(2'sd1),(2'd0)}?{((4'd0)?(-3'sd0):(2'd1))}:{((2'd0)?(4'd11):(4'sd1))});
  localparam signed [3:0] p15 = (4'd2 * (~^(~|(4'd10))));
  localparam signed [4:0] p16 = ((((3'd0)<<(-4'sd0))>>>(-((3'sd1)>>(-5'sd6))))<=(((-2'sd1)^(2'sd0))!==((2'sd0)|(5'd4))));
  localparam signed [5:0] p17 = {1{(5'sd7)}};

  assign y0 = {1{(2'd1)}};
  assign y1 = ((^(a3!==a5))>=((p10>=p1)-(p9&&p7)));
  assign y2 = (((|(b4>>a4))>>{2{(~&b2)}})^~(~^({1{(a2>>b3)}}===(~&(~&b3)))));
  assign y3 = {(&(~&p7)),(~^(^p3))};
  assign y4 = ((-(2'sd1))>>>((+(p8!=p7))!=((4'sd2)<(p16&&p4))));
  assign y5 = ((~(b0*b2))===(-(b1==a2)));
  assign y6 = (!((!{2{{3{b3}}}})<<{1{(!((~&b1)>=(~|p2)))}}));
  assign y7 = (!$unsigned((5'd2)));
  assign y8 = $unsigned({2{$signed($signed({{a5,b2,a0}}))}});
  assign y9 = {1{{1{(~((^b5)<<{4{b2}}))}}}};
  assign y10 = (+{b3,p1});
  assign y11 = {(4'd5),(3'd4),((p11<<<p16)<=(-2'sd0))};
  assign y12 = (+((!{((a4?a3:p10)?(b0?b3:p15):(b2<<<p4))})^{(~|b5),(|a0),(b2?b5:b4)}));
  assign y13 = ((2'd0)+(a5^a4));
  assign y14 = (-4'sd4);
  assign y15 = ($unsigned(((b0!==b1)))>(~^(~$signed((a2==a0)))));
  assign y16 = ((-(b4>>>a0))*(b5*b5));
  assign y17 = ((~{3{(p1>=p10)}})<<<{3{(~|(~^a3))}});
endmodule
