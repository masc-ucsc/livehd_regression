module expression_00625(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((3'd6)>(-3'sd3))};
  localparam [4:0] p1 = (-5'sd1);
  localparam [5:0] p2 = (~|{1{{1{(~{{4{(5'sd14)}}})}}}});
  localparam signed [3:0] p3 = ((~|((-4'sd0)?(5'd16):(3'd4)))?({(2'd2),(4'd11)}?(&(4'd10)):((4'd1)|(5'd14))):{((4'sd4)==(5'd1)),((2'd0)?(4'd0):(5'sd14)),{(4'sd3)}});
  localparam signed [4:0] p4 = (3'd1);
  localparam signed [5:0] p5 = ((((3'sd2)?(-4'sd6):(3'sd2))|((2'sd1)?(2'd1):(3'd1)))!=((((3'sd1)>>(-4'sd0))+(~(5'd20)))>>((4'd5)|((2'd2)^(3'd5)))));
  localparam [3:0] p6 = (-5'sd13);
  localparam [4:0] p7 = (((((2'sd0)>>(3'sd3))>((4'd14)/(4'd3)))==(((3'd6)^(2'd2))^~((-3'sd0)==(2'd3))))>>((((2'd3)<<(4'd12))+((-2'sd0)^~(5'd14)))<(((4'd2)==(-5'sd4))>>((2'd1)<=(5'sd9)))));
  localparam [5:0] p8 = (5'd11);
  localparam signed [3:0] p9 = ((+((4'd3)&(4'd8)))>=(+{3{(4'd13)}}));
  localparam signed [4:0] p10 = (((4'sd2)?(2'd1):(2'sd0))?((-5'sd8)?(3'sd2):(4'sd6)):{(5'd2 * (4'd8))});
  localparam signed [5:0] p11 = ((4'd14)?(-2'sd0):(5'sd8));
  localparam [3:0] p12 = ((5'd9)?(5'd22):(5'd3));
  localparam [4:0] p13 = (-((3'sd0)|(-3'sd0)));
  localparam [5:0] p14 = {1{(4'd3)}};
  localparam signed [3:0] p15 = {2{((~^(2'd3))-((-4'sd6)?(-2'sd0):(4'd14)))}};
  localparam signed [4:0] p16 = {1{{3{{(~|{(4'd3),(-2'sd0),(2'd2)})}}}}};
  localparam signed [5:0] p17 = ((4'd6)>(3'd7));

  assign y0 = ((((b1^p9)||(b0+p5)))<<<((5'd2 * (p14|p7))>=((+b3)||(a4))));
  assign y1 = ((+(((-a0)+$signed(a5))>>($unsigned((p12<<a1)))))^~(|((-((a2!=a4)/p11)))));
  assign y2 = {4{{1{(!(a1>>a1))}}}};
  assign y3 = $unsigned(({2{(b4!==b2)}}));
  assign y4 = (&((!((&a1)?(!a5):{2{b5}}))!=(-((+b1)&(-b5)))));
  assign y5 = (^{3{$signed((a1?b2:b3))}});
  assign y6 = ((p9<p13)?(p5>=p5):(p8?p11:p17));
  assign y7 = ((a4!==b2)>(3'd6));
  assign y8 = (({a0,a5}?{a0,a5,b0}:{p17,a5})=={3{{4{b1}}}});
  assign y9 = (|(~^(b2?b4:b2)));
  assign y10 = ({b5,a2,a1}!==(a5||b1));
  assign y11 = ((~&(&(b2?b0:b4)))!=(!(~^{4{b4}})));
  assign y12 = (($signed(a4)>>>$signed(b1))==={(~(a0|a3))});
  assign y13 = ({({b1}<={b3,a5})}==({a0,b3}||(b5&&a0)));
  assign y14 = $signed($signed({{(3'd3),(p4>>p10)},(3'sd2),($unsigned({p4,p0})>={p5,p16})}));
  assign y15 = {((5'd12)>($unsigned((-2'sd1))<={(b1?b5:p2)}))};
  assign y16 = ((~{(3'sd3)})?(5'd11):{(4'd8),$signed(a4),(b4?b4:b2)});
  assign y17 = (&{3{{2{p16}}}});
endmodule
