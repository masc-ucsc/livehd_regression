module expression_00336(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(|({(4'd0)}^(2'd3))));
  localparam [4:0] p1 = (-5'sd7);
  localparam [5:0] p2 = (((5'd12)==(3'd0))<<<(3'd1));
  localparam signed [3:0] p3 = ((&((5'd6)==(-4'sd4)))!==((5'd18)>=(-5'sd0)));
  localparam signed [4:0] p4 = ((3'sd1)<<<(3'd0));
  localparam signed [5:0] p5 = (~(((~|(|(4'd7)))>>((3'd5)<<<(5'd21)))==((~(&(5'd1)))<<((2'd0)===(5'sd8)))));
  localparam [3:0] p6 = (((-2'sd0)*((2'sd0)&&(5'd10)))<<<(((5'sd2)!=(-4'sd5))+(-4'sd1)));
  localparam [4:0] p7 = ((-((4'd0)?(4'd12):(4'd8)))?(((5'd30)?(-4'sd1):(-3'sd1))?((-5'sd9)?(-4'sd2):(4'd13)):((3'd6)?(-4'sd3):(4'd7))):(((3'd2)?(4'd8):(5'd16))?(-(3'd4)):(-(5'd0))));
  localparam [5:0] p8 = ((5'sd7)-(((5'd3)&&(3'sd3))>((4'd6)?(5'd13):(-4'sd4))));
  localparam signed [3:0] p9 = {{3{(5'd6)}},{(3'd0),(-4'sd6),(2'd1)}};
  localparam signed [4:0] p10 = (((-2'sd0)!==((2'd2)<<(5'sd4)))&(((3'd2)<=(4'sd2))==((2'd0)&(5'd12))));
  localparam signed [5:0] p11 = (~(-{({(2'd0)}<<((3'd2)?(5'sd4):(-3'sd1))),((~|(3'd1))&&((-4'sd4)<=(3'd3))),(((5'd2)?(2'sd0):(2'd0))===(~|(4'd3)))}));
  localparam [3:0] p12 = {{{{(2'd3),(5'd2),(-4'sd5)}},{3{(4'd11)}},{(-4'sd2),(3'd0),(3'd2)}}};
  localparam [4:0] p13 = {(2'sd0),(4'sd5),(-2'sd0)};
  localparam [5:0] p14 = ({((-3'sd2)^~(2'sd1)),((4'd12)?(-3'sd1):(2'd3)),(!(-3'sd0))}==({(4'd14),(5'd14)}|((-4'sd3)>(3'sd2))));
  localparam signed [3:0] p15 = (({3{(5'd20)}}?((4'd13)?(3'sd0):(5'sd7)):{(3'sd0)})&&(((5'sd14)==(3'd2))?((4'd14)?(2'd0):(-4'sd6)):(4'd2 * (5'd13))));
  localparam signed [4:0] p16 = ((~&(((2'sd1)==(3'd7))<<<(|(3'd4))))<=((~^(2'd3))*(~(-3'sd2))));
  localparam signed [5:0] p17 = {4{((3'd0)?(2'sd1):(-4'sd7))}};

  assign y0 = (5'd0);
  assign y1 = $signed(b1);
  assign y2 = ((~&((p10?a0:p11)?(-b0):(a4<p10)))?((~(&p1))<(p4?p9:p1)):(+((p1&&p11)-(~^b4))));
  assign y3 = ((2'd0)<(p10?b3:a2));
  assign y4 = $signed((b3!==a3));
  assign y5 = ((p11/p11)/p8);
  assign y6 = (6'd2 * (4'd14));
  assign y7 = (2'sd0);
  assign y8 = (2'd3);
  assign y9 = {(3'sd0),(a2?p7:a1)};
  assign y10 = ((-(~^(!$signed((b5?a3:b2)))))?((p7>>>a0)?(~|a2):(3'd3)):((~p0)?(p8?p8:b3):(p3?b0:p4)));
  assign y11 = {p11,p15,p0};
  assign y12 = {(-(((+(p4>=p3))>>(~(p8<a3)))>>>(-{$unsigned((&a3)),(p4>>a5),$signed((p15<p7))})))};
  assign y13 = {((p7<=p3)<<<(~b0)),((^a5)==={a3,b2,a1})};
  assign y14 = ((|$unsigned(p10))<(~^(p15|p11)));
  assign y15 = {4{(a4!==b3)}};
  assign y16 = {(-(|(~&(~|(~&p0))))),({p10,a2}?(!b4):(p11^p15))};
  assign y17 = ((2'sd0));
endmodule
