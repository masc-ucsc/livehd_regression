module expression_00235(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{2{(2'd2)}},{2{(5'd13)}},((5'sd7)^~(-3'sd2))};
  localparam [4:0] p1 = ((2'd2)?((3'sd2)?(4'd0):(5'sd4)):{(3'd6),(3'd7)});
  localparam [5:0] p2 = {{(5'sd4),(5'd27)},((2'd3)!==(5'd5)),((-2'sd0)>>>(-4'sd3))};
  localparam signed [3:0] p3 = ({(-2'sd1),(5'd22),(2'sd0)}?{2{((5'd23)?(4'd6):(-4'sd6))}}:(5'd2 * ((3'd5)?(4'd5):(5'd4))));
  localparam signed [4:0] p4 = {(({3{(5'd0)}}^{4{(-5'sd10)}})<(-(~&{4{(5'sd6)}})))};
  localparam signed [5:0] p5 = {1{(4'd5)}};
  localparam [3:0] p6 = (^(((4'd9)?(2'sd1):(-4'sd7))?(~|(4'd13)):(~&(3'd3))));
  localparam [4:0] p7 = ({(6'd2 * (5'd16))}-((+((5'd26)&(2'd3)))===(2'd2)));
  localparam [5:0] p8 = ((-5'sd12)!=(5'sd13));
  localparam signed [3:0] p9 = (&(5'd15));
  localparam signed [4:0] p10 = {4{(4'd6)}};
  localparam signed [5:0] p11 = {2{{{(2'd0),(5'd8)},{1{{3{(2'sd1)}}}},{(5'd31),(-5'sd11),(5'd8)}}}};
  localparam [3:0] p12 = (6'd2 * (2'd0));
  localparam [4:0] p13 = (-3'sd2);
  localparam [5:0] p14 = {2{{1{{((2'sd0)^(4'd9))}}}}};
  localparam signed [3:0] p15 = (({(2'd3),(-3'sd3),(2'd0)}>=(4'd2 * (5'd1)))|(~^((&((-4'sd4)<<<(3'd4)))<<<{(-5'sd13)})));
  localparam signed [4:0] p16 = ({(((2'sd1)-(2'sd0))-((-2'sd0)?(-5'sd10):(3'sd3)))}>>>({(-5'sd12),(4'd7),(-2'sd1)}?((2'sd0)!==(-3'sd1)):((4'sd7)?(3'd2):(4'sd2))));
  localparam signed [5:0] p17 = (~^{(+((-4'sd1)&(4'd8))),(!(~^(-5'sd4)))});

  assign y0 = (3'sd1);
  assign y1 = (p12^~p0);
  assign y2 = {4{a4}};
  assign y3 = ({2{$signed(b1)}}<=($signed(a0)<<{4{a3}}));
  assign y4 = ((^$unsigned((3'd4)))||(~^((3'd3)>>>($signed(b4)&&$signed(p13)))));
  assign y5 = {b1,b5};
  assign y6 = (((b4?b4:b0)===(a0>=a5))?((a0?b5:a2)<<<(b4?p10:p4)):((p10?a2:a0)%a3));
  assign y7 = ($signed(((-5'sd9)===$signed(((|a0)))))>>({(-5'sd3),{p0},(~|b2)}&&{(~&p11),(p0>p4)}));
  assign y8 = (((^(p9?b4:b1))/p15)+(((-p3)==(p12?b5:p12))^~(+(~&(-p6)))));
  assign y9 = (2'd0);
  assign y10 = {4{((&a2)?(-p0):{1{b3}})}};
  assign y11 = ((4'd1)!=(+b1));
  assign y12 = (5'd0);
  assign y13 = (p10^~p3);
  assign y14 = (5'd30);
  assign y15 = $unsigned($signed((-5'sd10)));
  assign y16 = (-(!{2{({2{a1}}?(a2?p7:b5):(&b4))}}));
  assign y17 = (((a1!==b2)==(a3!=p9))+({4{p14}}<=(a0<b5)));
endmodule
