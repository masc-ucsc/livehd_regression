module expression_00884(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'sd3)?(4'd3):(3'sd3))?(!(5'd14)):(&(5'd4)));
  localparam [4:0] p1 = (((5'sd8)||(-2'sd1))||(2'd1));
  localparam [5:0] p2 = ((((-5'sd10)?(5'd9):(-3'sd2))>=({4{(3'd0)}}<<<((3'd5)||(4'sd2))))-(&({2{(4'd12)}}?((5'd14)+(2'sd0)):{1{(-5'sd13)}})));
  localparam signed [3:0] p3 = (5'd2);
  localparam signed [4:0] p4 = (((4'd14)^(-5'sd5))?((3'sd1)?(2'd3):(4'd7)):((4'd13)>>(-5'sd7)));
  localparam signed [5:0] p5 = {(4'sd0),(2'sd0)};
  localparam [3:0] p6 = ({2{(4'd13)}}<<(2'd3));
  localparam [4:0] p7 = {(5'd20),(5'sd6)};
  localparam [5:0] p8 = (2'sd1);
  localparam signed [3:0] p9 = (+((6'd2 * ((2'd1)>>>(3'd5)))+(((5'd28)?(5'd19):(3'd0))?((4'd2)/(4'd11)):((-3'sd0)===(2'd0)))));
  localparam signed [4:0] p10 = ((-(|(-5'sd11)))/(3'sd3));
  localparam signed [5:0] p11 = {(((3'd7)-(5'd4))&((3'd5)||(2'sd0)))};
  localparam [3:0] p12 = (((2'sd0)?(5'd13):(4'd2))?(!((4'd5)==(3'd4))):(4'd2 * (4'd3)));
  localparam [4:0] p13 = ((-4'sd4)?(-5'sd7):(3'd7));
  localparam [5:0] p14 = (!(|(~&((~|(!(!(!((4'sd3)^~(-5'sd7))))))!==((~^(3'd4))?((2'd3)?(-2'sd0):(2'd0)):(^(-4'sd0)))))));
  localparam signed [3:0] p15 = {(3'd6)};
  localparam signed [4:0] p16 = {{4{(3'd3)}},{(((5'sd15)>(3'd1))||{(3'sd1),(5'd23),(2'sd1)})}};
  localparam signed [5:0] p17 = {(({{(-5'sd5),(2'sd0)}}&&{4{(3'd6)}})&(~^{(^{(4'sd3),(4'd5)})}))};

  assign y0 = ({(b5?a3:b1)}<<<(a1?b5:b2));
  assign y1 = (~&$signed({2{$unsigned((!(|(!$signed(p9)))))}}));
  assign y2 = (~&(4'd0));
  assign y3 = ((5'd2 * (a0<<<p0))&&$signed((-4'sd6)));
  assign y4 = {(5'd28)};
  assign y5 = (b3);
  assign y6 = (p2?p12:p8);
  assign y7 = ({{4{p12}}}?{(!{3{b3}})}:(-{b1,p5}));
  assign y8 = ((~(a2&&b4))<<<(p4==a0));
  assign y9 = (((-$signed((a5?p3:a3)))?{2{(a5)}}:{2{(a5<=b2)}}));
  assign y10 = (p11>>>p13);
  assign y11 = ((-(b3?b2:a0))!==(b5>=a0));
  assign y12 = ((b0?p15:p6)?((a5?a5:p8)):(p14?p15:p14));
  assign y13 = (~|{2{((^(b5^~b4))&&(a4>>>a0))}});
  assign y14 = ({4{{p14,p3,p16}}}<<<{{{(~|p0),(b0!==a0)},(4'd2 * {p7})}});
  assign y15 = ({{p7,b1,a1},$unsigned((a2))});
  assign y16 = {3{p9}};
  assign y17 = (|{1{({1{(3'sd0)}}<={{4{a5}},(a4+p8),(3'd3)})}});
endmodule
