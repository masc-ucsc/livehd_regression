module expression_00217(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((5'd29)?(3'd4):(-2'sd1))&&((-2'sd1)-(4'sd0)));
  localparam [4:0] p1 = (((2'd0)?(-4'sd3):(-4'sd1))?((3'd2)?(4'd11):(3'sd1)):((2'd1)?(2'sd1):(4'd7)));
  localparam [5:0] p2 = (((-4'sd4)|(3'd7))?((2'd1)!==(4'sd6)):(~&((-4'sd2)>>(4'd9))));
  localparam signed [3:0] p3 = {3{({(-4'sd2),(3'sd1)}?((5'sd1)?(4'd8):(5'd20)):((-3'sd1)?(2'd1):(-2'sd1)))}};
  localparam signed [4:0] p4 = (~(((-4'sd3)?(2'd1):(3'd3))?(((-4'sd7)<<<(4'd1))!=((2'sd0)&(5'd15))):{1{((4'sd0)?(4'sd5):(3'd4))}}));
  localparam signed [5:0] p5 = {2{({(4'd8),(2'd0)}&{(-4'sd4),(3'd4),(2'd1)})}};
  localparam [3:0] p6 = ((3'd3)?(4'd10):(5'd16));
  localparam [4:0] p7 = ((~|((-(3'd1))^{(2'sd0),(4'd14),(3'd0)}))|(((4'sd7)-(2'd0))^(&(3'd4))));
  localparam [5:0] p8 = (((4'd12)!=(-3'sd0))<={2{(2'sd0)}});
  localparam signed [3:0] p9 = (+{4{(2'd0)}});
  localparam signed [4:0] p10 = ((((3'sd3)===(3'd0))==(~&(2'd3)))>((3'sd0)?(5'd1):(3'sd1)));
  localparam signed [5:0] p11 = ((((-4'sd1)<(2'sd0))^~((5'd14)>(-4'sd7)))<<{((-5'sd11)<=(-2'sd0)),((5'd14)||(-3'sd3))});
  localparam [3:0] p12 = {(2'd1),(-5'sd15),(3'sd2)};
  localparam [4:0] p13 = ((^(~^((3'sd1)!=(-5'sd7))))?(~((5'd10)?(3'd3):(2'd2))):(~(|((3'd7)!=(4'd0)))));
  localparam [5:0] p14 = {3{{1{{(-2'sd0),(4'd3),(-3'sd0)}}}}};
  localparam signed [3:0] p15 = {{({(4'd4)}<{(5'd0),(5'd28)})},({1{(5'd29)}}?((4'd2)^(-5'sd14)):((5'd22)!==(5'd3)))};
  localparam signed [4:0] p16 = (3'd3);
  localparam signed [5:0] p17 = ((5'd29)||(4'sd3));

  assign y0 = (p11?p13:b2);
  assign y1 = {4{{{2{p16}}}}};
  assign y2 = (((b1*b3)?(~^a2):(b0?b3:p16))&(~|((&a0)?(b3?p5:b3):(-b4))));
  assign y3 = (p12^~p7);
  assign y4 = ({2{b0}}!={2{p15}});
  assign y5 = (((b5<<a5)/b4)+((4'd2 * p14)/b2));
  assign y6 = ((5'd6)>>((a3?p16:a1)==(4'd10)));
  assign y7 = (2'sd1);
  assign y8 = (2'd0);
  assign y9 = ({b1,p9,p5}^~(4'd10));
  assign y10 = ((a3&b0)<=(a3<=b0));
  assign y11 = {4{(b5?a2:a1)}};
  assign y12 = (((-p13)^~(-5'sd6))<<({b2,p5,p14}^(5'sd4)));
  assign y13 = {3{(a1?p10:b5)}};
  assign y14 = ({({b3,a2}),$signed($signed(a2))}?(($unsigned(p15)?(a1?b0:p13):{p0})):{$unsigned(p17),(b4?b3:b4),(b0)});
  assign y15 = {2{({b0}^~{1{b3}})}};
  assign y16 = (&p16);
  assign y17 = {a3,p3,p0};
endmodule
