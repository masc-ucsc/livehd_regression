module expression_00099(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-3'sd2)?(-2'sd1):{((4'sd2)!==(5'sd7))});
  localparam [4:0] p1 = (~^(-5'sd0));
  localparam [5:0] p2 = (+{((2'd1)>(-3'sd0)),(+(4'd12)),{(3'd5)}});
  localparam signed [3:0] p3 = (((4'd6)?(-5'sd2):(5'd17))?({(5'sd11),(4'd4),(5'sd10)}<<<((-2'sd1)?(3'sd2):(2'd1))):({(3'd1),(-2'sd0)}<={(-2'sd0)}));
  localparam signed [4:0] p4 = (|((~^(5'sd4))^(~|(-5'sd13))));
  localparam signed [5:0] p5 = (~^(~{{(4'sd2),(2'd1)}}));
  localparam [3:0] p6 = (4'd2 * (3'd0));
  localparam [4:0] p7 = ((~^{(2'd3),(2'd1),(-2'sd1)})?(~&(~|(3'd7))):{(3'sd1),(4'd12),(-4'sd6)});
  localparam [5:0] p8 = (-5'sd0);
  localparam signed [3:0] p9 = ((-3'sd2)!=(5'd24));
  localparam signed [4:0] p10 = ((4'd2 * ((3'd5)==(3'd3)))?(((-2'sd1)|(2'd1))?{(2'd3),(3'd0)}:{1{(5'd8)}}):(!{((2'sd0)<<<(-4'sd1)),{(2'sd0)}}));
  localparam signed [5:0] p11 = (((4'd6)<(2'd1))-(!(-4'sd4)));
  localparam [3:0] p12 = (((3'd4)<(3'sd3))>=((4'sd1)+(5'd1)));
  localparam [4:0] p13 = ({{{(5'd15),(3'sd2),(-5'sd2)}}}?((3'd4)?(5'd20):(3'd4)):(((3'd5)?(-4'sd7):(2'd2))^~{(2'd0),(3'sd1),(4'sd7)}));
  localparam [5:0] p14 = ((|(-3'sd3))!=((-2'sd1)===(3'd0)));
  localparam signed [3:0] p15 = (6'd2 * ((4'd15)|(4'd13)));
  localparam signed [4:0] p16 = {2{((4'd7)?(-4'sd4):(2'sd1))}};
  localparam signed [5:0] p17 = (((5'd13)^{(2'sd1),(-3'sd3),(-5'sd8)})^~(6'd2 * ((2'd0)>>(4'd9))));

  assign y0 = ((+b3)-{p7,a3,p13});
  assign y1 = ((a0-b1)^~(b5?b4:a1));
  assign y2 = {2{(2'sd0)}};
  assign y3 = (p1?p13:p2);
  assign y4 = {4{b1}};
  assign y5 = ({(a2&b2),(a2===b5),(a4!==b1)}==(!({(3'sd3)}?{a2,b4}:(a0>b0))));
  assign y6 = (6'd2 * {{b0,b1,a1}});
  assign y7 = {4{({4{a3}})}};
  assign y8 = (4'sd6);
  assign y9 = (4'sd7);
  assign y10 = ((((b5||a1)>>>(a5<=a4))||(b0?b0:b2))^~{(~^(b2?a5:b5)),(p5<<b4),(b5?b3:b1)});
  assign y11 = ((^(+((b3<<<p0)>>>(p14&p10))))^~(|((a5==p4)!=(b0!==a3))));
  assign y12 = ({$signed((~&(~^(&(~&{p0})))))});
  assign y13 = ((p12^p6)?(p0?b5:p12):(p0));
  assign y14 = (((2'sd0)?(p15!=b0):(p2?a3:p7))&&(-2'sd1));
  assign y15 = (~|(((p6^p1)==(~|{1{p3}}))^~({1{p9}}?{2{p10}}:(p4==p1))));
  assign y16 = {3{({2{p7}}>>(5'd30))}};
  assign y17 = (p11^~p3);
endmodule
