module expression_00741(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(~^((|(~|(~&(-2'sd1))))?{((4'sd0)?(2'd3):(5'd13))}:{1{((5'd24)&&(5'd14))}})));
  localparam [4:0] p1 = (~(((~^(-4'sd4))^((3'd5)!=(5'sd15)))+((|(2'd0))+((5'sd8)===(3'd0)))));
  localparam [5:0] p2 = (-(~((3'd5)&(-4'sd4))));
  localparam signed [3:0] p3 = (((3'sd0)?(5'd27):(-3'sd1))?((5'd13)?(-3'sd1):(2'd1)):((5'd1)?(3'd0):(2'd2)));
  localparam signed [4:0] p4 = (4'd9);
  localparam signed [5:0] p5 = (({(5'sd1),(3'd4),(2'd0)}!==(|(4'sd5)))>>({1{(4'd8)}}&((2'd0)<<<(2'sd0))));
  localparam [3:0] p6 = {{(5'd11),(2'd2),(2'sd1)},((5'sd0)!=(-5'sd10)),((-4'sd5)<<(2'd3))};
  localparam [4:0] p7 = (((!(4'sd5))?((4'sd0)==(-5'sd13)):(~^(-3'sd3)))<(((4'd13)?(2'd1):(2'd2))!=((-3'sd0)!==(2'd0))));
  localparam [5:0] p8 = ({(~&(-4'sd1))}&&((4'sd3)?(4'sd5):(3'sd3)));
  localparam signed [3:0] p9 = ((-2'sd1)==(-4'sd2));
  localparam signed [4:0] p10 = (5'd8);
  localparam signed [5:0] p11 = (3'sd3);
  localparam [3:0] p12 = ((~|(|(~|(4'sd4))))?(((2'sd1)?(-3'sd0):(-5'sd15))-{2{(-4'sd7)}}):{(3'sd1),(3'd1),(4'sd4)});
  localparam [4:0] p13 = ((((2'd2)>(4'd14))^~((4'd2)||(4'd0)))>>>{{((-5'sd6)>>(5'sd2)),{(3'sd1)}}});
  localparam [5:0] p14 = ((-(3'd0))?{(3'sd3),(5'sd7)}:((-5'sd8)|(3'sd0)));
  localparam signed [3:0] p15 = (~|(((2'sd1)-(2'sd1))+((5'sd12)==(3'd5))));
  localparam signed [4:0] p16 = {2{{3{(5'd19)}}}};
  localparam signed [5:0] p17 = (+(|(~|{{4{{(~^(5'sd9))}}}})));

  assign y0 = (-4'sd0);
  assign y1 = (({a3,p6}?(|b3):(-b0))?(-{(-p9),(b0<<<b0),{p13,a1}}):(^({p16}?(+p16):(~p11))));
  assign y2 = (a2*p17);
  assign y3 = ((^a1)?$signed(p2):(+b0));
  assign y4 = (6'd2 * {a2,p13,a0});
  assign y5 = ((-3'sd0)?(a4===b3):(p14?p9:p5));
  assign y6 = $unsigned($unsigned((p13?p11:p0)));
  assign y7 = {({4{a5}}!=={(a0&b4),(+a4)})};
  assign y8 = (|(~&((-(~&((b0/a3)>(a0>>>b0))))||(((p0<<a2)>>>(p12&b4))^((b2>>>a3)===(b3<a1))))));
  assign y9 = $signed((($unsigned((-a4))<<(a4<=b1))^~((a4>a2)>(6'd2 * b2))));
  assign y10 = ({(^({(b4!==b1)}|(a2?p1:a3)))}>((a4===a1)?(b1||b2):(-(+p14))));
  assign y11 = {((a5?a2:b1)?(b0?b3:b2):(~^a4)),{(~(4'd5))}};
  assign y12 = {{((p3?p7:p8)?(b0?b4:p6):{(|a5)}),((~|(p2?p5:p15))?(~^(p9?b0:p17)):{p11,b0})}};
  assign y13 = (~|(&{3{((3'd5)^(a4>>a1))}}));
  assign y14 = ((-3'sd2)?(~&{p17,p12,p16}):{(p13?p7:p8)});
  assign y15 = (2'd2);
  assign y16 = (((^(-3'sd1))&(+(+(~b5))))!==(~|(+(!(~(~&(^(~b1))))))));
  assign y17 = {2{(-{3{(-p12)}})}};
endmodule
