module expression_00742(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!{(|((4'd13)!=(4'd11))),(&(-((3'sd1)<(4'd8)))),(~(~&(~&(5'sd5))))});
  localparam [4:0] p1 = ((5'd6)^((5'd17)<=(5'd16)));
  localparam [5:0] p2 = ({4{(5'd2)}}?{1{(3'd5)}}:((2'sd1)?(2'd3):(2'd2)));
  localparam signed [3:0] p3 = {((2'sd0)>=(3'sd3)),{(4'd0),(2'sd1),(5'd8)}};
  localparam signed [4:0] p4 = ((5'sd11)<<(3'sd2));
  localparam signed [5:0] p5 = ((4'd5)?(4'sd4):(-5'sd6));
  localparam [3:0] p6 = {{((-3'sd3)?(4'sd3):(-5'sd11))}};
  localparam [4:0] p7 = ({(3'd6),(5'd6),(2'd1)}!=(|(~^(5'd12))));
  localparam [5:0] p8 = ((((4'd0)?(2'sd1):(2'd3))<<(+{3{(5'd7)}}))&{3{(-(-5'sd7))}});
  localparam signed [3:0] p9 = ((5'd2 * (3'd5))<<((-3'sd2)<=(3'sd2)));
  localparam signed [4:0] p10 = {{(4'd14),(4'sd4),(4'd6)}};
  localparam signed [5:0] p11 = {(~&{(-(~(2'd2))),(|{(4'sd2)})}),(~^(~{(+(4'sd4)),(!(5'd7)),(~|(-5'sd15))}))};
  localparam [3:0] p12 = (2'd3);
  localparam [4:0] p13 = (&{(4'd14),(-3'sd3)});
  localparam [5:0] p14 = ({((5'd22)?(3'd5):(4'd15)),{(-3'sd2),(-4'sd4),(-2'sd1)}}==({(3'd6)}?((5'd2)>>(2'sd0)):((5'd13)>>>(3'd4))));
  localparam signed [3:0] p15 = ((5'd23)?(5'd10):(4'sd7));
  localparam signed [4:0] p16 = {2{(5'd5)}};
  localparam signed [5:0] p17 = (!((4'd3)&(4'sd3)));

  assign y0 = (~|$signed(($unsigned(((b2===b2)))&((p3<<<p6)>>>{3{b1}}))));
  assign y1 = $signed($unsigned((~&a0)));
  assign y2 = {(~^((p12+b5)<<<(p10||p5)))};
  assign y3 = (3'd1);
  assign y4 = (|({{4{p8}},(p9?b2:b4),(b4>>>p3)}==(^{2{({a1}+(p0?p5:p13))}})));
  assign y5 = (~{4{p3}});
  assign y6 = ((p8?b2:b4)?(p7?b1:b4):{p1,b0,p5});
  assign y7 = (a4===a5);
  assign y8 = (~&(4'd12));
  assign y9 = ((+((p14||p16)<=(~|(5'd22))))&(&{4{(!p5)}}));
  assign y10 = (5'sd8);
  assign y11 = (~^((~((p8>>b4)-(~^{p15,p4})))>>>{(p11>=p6),(+(p12^~p14))}));
  assign y12 = (5'd9);
  assign y13 = {(-(~^((p15^~p5)>=(|a0))))};
  assign y14 = (~|(&(|{1{(~|((-({3{a1}}))==(-(^{2{p2}}))))}})));
  assign y15 = {b3,b2,b5};
  assign y16 = {4{a2}};
  assign y17 = (^(~|(~((~&(~&a5))?(-(!b4)):(^(^b0))))));
endmodule
