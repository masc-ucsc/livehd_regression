module expression_00072(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'd8);
  localparam [4:0] p1 = (!(!(2'sd1)));
  localparam [5:0] p2 = {4{{2{(2'sd0)}}}};
  localparam signed [3:0] p3 = ((5'd30)&(5'd7));
  localparam signed [4:0] p4 = (~^(+{(3'd4),(-2'sd1),(4'sd3)}));
  localparam signed [5:0] p5 = {(&(~(-((2'd0)<(2'd2)))))};
  localparam [3:0] p6 = ((((4'd5)?(4'd10):(4'sd7))^(6'd2 * (3'd3)))!=={((4'sd7)?(5'd28):(4'd4)),((4'd14)?(-3'sd0):(4'd15))});
  localparam [4:0] p7 = {1{(-4'sd2)}};
  localparam [5:0] p8 = (5'sd12);
  localparam signed [3:0] p9 = (2'd1);
  localparam signed [4:0] p10 = (~(~&(+(4'd10))));
  localparam signed [5:0] p11 = (~&(3'd0));
  localparam [3:0] p12 = {(-(2'sd1))};
  localparam [4:0] p13 = (((-3'sd0)?(2'd1):(3'd2))?{(-5'sd6)}:{(2'd1),(4'd9),(-3'sd0)});
  localparam [5:0] p14 = (((~^(2'sd0))?((4'd0)>>(3'd0)):(3'sd0))^(~|(4'sd4)));
  localparam signed [3:0] p15 = (|(!(+((((-4'sd1)/(4'd15))==(~^(4'd4)))&&(!((&(2'd2))+((3'sd2)||(3'd5))))))));
  localparam signed [4:0] p16 = (~&(-2'sd1));
  localparam signed [5:0] p17 = {(~|(((4'sd7)>>>(5'sd12))<=(+{(-2'sd1),(2'd1),(5'd10)}))),({(3'sd3),(4'sd3),(4'd6)}|(&(~&(~^(4'd13)))))};

  assign y0 = ((a4<p12)<<(p13-b3));
  assign y1 = ((&({2{p4}}?(p10?p1:p10):(p13?p5:p12)))?(&{2{(|p12)}}):(&{4{p3}}));
  assign y2 = ({4{b3}}<={1{(!(a4===a1))}});
  assign y3 = ((2'd2)?(5'd2 * (~(^b2))):({a4,b4}>=(b2?a3:a1)));
  assign y4 = (+(!{4{(!(~&{p1}))}}));
  assign y5 = (((b4?p3:b0)?(p16?p3:p11):(a5?b1:b2))?((a3?a3:b2)?(b4?p3:p2):(b0?b4:a0)):((a3?p7:p4)?(a0?p1:p2):(p2?p16:p1)));
  assign y6 = (5'd12);
  assign y7 = (b2>>a1);
  assign y8 = (&(~|(^(-(~p17)))));
  assign y9 = (~($signed((&(b5==a1)))<=((a5)>=$unsigned(a3))));
  assign y10 = ((3'sd2));
  assign y11 = {{{b3,b3},{p13,b3,a0},{p7,p6}},{{{p0,b2},{p0}},{p4,p15,b0}}};
  assign y12 = ((|(~^((b5&b5)/p1)))>((~|(a5<<b2))!==(!(b3*b5))));
  assign y13 = (~(((~b3)/a1)<<<((|p17)-(p6>>>p1))));
  assign y14 = (^{{p10,p5,p13},((!p12)!=(p9^p5)),(~|{b1,p14,p10})});
  assign y15 = (|(~|(((p8||b5)?(&(~|p9)):(p9==a2))>={3{{1{(p15-p16)}}}})));
  assign y16 = (~&(-(~(&(^(~^p6))))));
  assign y17 = (p8?a5:p9);
endmodule
