module expression_00980(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(!(5'd18)),((4'd2)==(2'd0)),{3{(-3'sd3)}}}};
  localparam [4:0] p1 = (-3'sd2);
  localparam [5:0] p2 = (|(5'sd12));
  localparam signed [3:0] p3 = (~((~^(!(3'sd3)))?(-(!(-2'sd0))):(~&((2'sd0)?(2'd2):(2'sd1)))));
  localparam signed [4:0] p4 = (-((!((-5'sd6)?(2'sd0):(3'sd2)))?{3{(3'sd3)}}:{2{(-2'sd1)}}));
  localparam signed [5:0] p5 = (~((5'd22)>>>{4{(-3'sd2)}}));
  localparam [3:0] p6 = (5'sd9);
  localparam [4:0] p7 = {{(-3'sd0),(3'd1)}};
  localparam [5:0] p8 = (-(2'd2));
  localparam signed [3:0] p9 = {1{(4'd9)}};
  localparam signed [4:0] p10 = (-2'sd1);
  localparam signed [5:0] p11 = {(3'd3),(4'd5)};
  localparam [3:0] p12 = {3{(4'sd1)}};
  localparam [4:0] p13 = (((2'd2)&((2'sd1)<<<(5'd14)))!=(!(!(5'sd15))));
  localparam [5:0] p14 = {(((-3'sd2)>>>(3'd1))!=((3'sd1)?(-5'sd4):(3'd0))),(((5'd23)&(-3'sd0))^(&(5'd14))),(((3'd7)<<(2'sd1))>>>{(2'd1),(5'd30)})};
  localparam signed [3:0] p15 = {1{((-3'sd1)+(3'sd1))}};
  localparam signed [4:0] p16 = (+{(+(^(2'd3))),{1{{(5'd13),(-5'sd8)}}},{3{(5'sd0)}}});
  localparam signed [5:0] p17 = (((4'd15)^(2'd3))|(^((3'd2)?(5'd15):(3'sd1))));

  assign y0 = ((~|(~(~(&(!(~&(!(p13?p7:p7))))))))|(~&(&(~&((+p7)?(a0<<<p6):(p5?p4:p7))))));
  assign y1 = ($unsigned((!p16))^(p15-p4));
  assign y2 = ($signed(p13)<<<{p17,b3,b2});
  assign y3 = ((&(~{b5,b2,p10}))>>>((b1==a2)!=={(&a1)}));
  assign y4 = (5'd2 * (^(~|a2)));
  assign y5 = (($unsigned($unsigned(($unsigned(b4)&&(b2>b3))))!==$signed(($unsigned((4'd2 * b1))+((a1^b3))))));
  assign y6 = {2{{3{a5}}}};
  assign y7 = (a2===a5);
  assign y8 = ((5'd0)^((~&(4'd2 * b2))!=(4'sd3)));
  assign y9 = (~|(3'sd0));
  assign y10 = (b0^~b5);
  assign y11 = (((a0>>p10)>(p17?b1:p2))>>{3{{4{p13}}}});
  assign y12 = $unsigned((~|(~&(!({4{a5}}>>>(a5))))));
  assign y13 = {3{(4'd6)}};
  assign y14 = ((($signed((p14&p12))&$unsigned((p5)))?($signed((a3>>b3))^~(p9<<<b5)):((p5?p11:p13)%p7)));
  assign y15 = {((a4?b4:p7)>(p10?b4:p17)),((p1>=p2)!=(b1===a4)),{((p2==a2)<=(p0|a1))}};
  assign y16 = (((4'd5)||(b3<=p6))>>(a0?a4:a1));
  assign y17 = (p12>>>p17);
endmodule
