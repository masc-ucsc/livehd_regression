module expression_00245(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(~(+(((3'sd3)>>(-5'sd11))>(!((3'd2)?(5'd22):(-2'sd0)))))),(+((-{(-3'sd2),(4'd2),(3'd6)})||(+((5'd4)^(5'd3)))))};
  localparam [4:0] p1 = ((^(((4'sd2)-(3'sd1))?((5'd24)<=(4'd10)):(~|(-3'sd2))))<=(-((^(3'sd1))?((3'sd0)<<<(5'd27)):((4'sd0)!==(-2'sd0)))));
  localparam [5:0] p2 = (-2'sd0);
  localparam signed [3:0] p3 = (5'd2 * (4'd12));
  localparam signed [4:0] p4 = ((3'd7)?(2'sd1):(3'sd2));
  localparam signed [5:0] p5 = ((~&(~(~|(2'sd0))))?(4'd3):(~|(4'd2)));
  localparam [3:0] p6 = ((^(~(~(4'd15))))?(((2'd3)?(3'd5):(4'sd0))>>(^(5'sd11))):((|(-5'sd1))-((4'd2)+(2'sd1))));
  localparam [4:0] p7 = {1{(4'sd0)}};
  localparam [5:0] p8 = (((~&{{(2'd2),(4'sd7),(-2'sd0)}})>>>(((5'd3)===(2'd3))<={(2'd3),(5'd3)}))+{(((2'd0)&&(-2'sd0))?{(3'd5),(-3'sd2)}:(~|(3'd7)))});
  localparam signed [3:0] p9 = {4{{4{(-2'sd0)}}}};
  localparam signed [4:0] p10 = (~|((-3'sd2)&(-(~^(^(2'd0))))));
  localparam signed [5:0] p11 = {4{{1{((2'd0)||(4'sd5))}}}};
  localparam [3:0] p12 = {({(4'd10)}^~(-2'sd1)),{{(5'd19),(5'd6)}},{{(-5'sd13),(2'd3)},((-3'sd1)|(3'd2))}};
  localparam [4:0] p13 = {((2'sd0)<(~|(-3'sd3)))};
  localparam [5:0] p14 = (((2'd0)===(5'd5))+((-4'sd0)!==(2'd2)));
  localparam signed [3:0] p15 = (~&(!(+(&(&(!(+(!(+(~(^(~|(~(!(+(2'sd0))))))))))))))));
  localparam signed [4:0] p16 = ((4'sd5)|(2'd3));
  localparam signed [5:0] p17 = {(4'd5),(4'sd2),(4'd15)};

  assign y0 = ((4'sd3)-((5'd18)<(~&(4'sd6))));
  assign y1 = ((&(~^(|$signed({3{(2'sd1)}})))));
  assign y2 = ((((b5>=b4)<<{b1,a1,a1})-$unsigned({b5,a1,a0}))===({(b0),(a0<=a2)}+{(a4>>>b2),$unsigned(a4)}));
  assign y3 = ({2{p6}}>(a0+p13));
  assign y4 = ((~^b4)==={a3});
  assign y5 = {({2{({4{b4}}===$signed(b5))}}<<<({{{p9}}}!=((b5<<<p0))))};
  assign y6 = {3{(4'd5)}};
  assign y7 = (5'd2 * $unsigned((p13?a5:a4)));
  assign y8 = ((((&b5)?(a4?b2:a3):(~p7))||((a3>p2)?(b0^~p14):(p13>>>p11)))&(((b1?b2:a2)^(a2||b3))+((a1+a2)?(p3==b4):(p11?p11:p5))));
  assign y9 = (4'd5);
  assign y10 = (((4'd1)?(p15?p14:p12):(b4<<p1))?$unsigned($unsigned((p7?p6:p15))):(!((~&b2)!=(p6+p4))));
  assign y11 = (~|(b1!==a3));
  assign y12 = ((b2?b0:p10)?{p6}:(2'sd0));
  assign y13 = $unsigned({2{{(&p2)}}});
  assign y14 = (+(p3-p1));
  assign y15 = ((-{a0,a1,a4})?(~^{p10,p0,a2}):{(&b4),(p12==b5)});
  assign y16 = (~(-(+$unsigned($signed((-3'sd0))))));
  assign y17 = (-$unsigned((-(^(({p12}?(~^b1):(|p13))?({p14,p5}?(!p1):$signed(p9)):$signed((|{p12,p8})))))));
endmodule
