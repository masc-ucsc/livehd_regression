module expression_00693(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd1)?(5'sd8):(3'd5))<=(~|(|(5'd11))));
  localparam [4:0] p1 = {2{(2'd0)}};
  localparam [5:0] p2 = {((4'd12)===(2'sd1)),{(5'd21),(3'sd1)},((3'd1)&(-2'sd0))};
  localparam signed [3:0] p3 = ((((~&(3'sd0))<=(-4'sd2))&&{1{(3'sd0)}})^~({1{{3{(3'd0)}}}}>=(-5'sd8)));
  localparam signed [4:0] p4 = (|((|(~(5'd2)))?((2'sd0)?(-3'sd1):(2'd3)):(^((2'sd1)?(2'd2):(2'd3)))));
  localparam signed [5:0] p5 = (5'd2 * ((3'd2)&&(5'd29)));
  localparam [3:0] p6 = (&((-2'sd1)?(4'd12):(5'd28)));
  localparam [4:0] p7 = ((((-4'sd6)^~(-5'sd4))?((4'd15)^~(4'sd4)):((2'd2)?(2'd3):(4'd5)))?(((-5'sd8)==(4'd2))?((3'd5)>>>(3'd7)):((2'sd1)?(2'sd1):(4'sd7))):(((5'sd14)|(3'sd2))?((-2'sd1)?(2'sd1):(4'd4)):((2'sd0)?(-5'sd7):(5'd16))));
  localparam [5:0] p8 = (+{4{((3'sd3)^(4'd4))}});
  localparam signed [3:0] p9 = {(((4'd13)?(4'sd0):(5'd0))==((5'd18)>>(-2'sd0))),(((3'd5)<=(-3'sd2))||((5'd16)||(3'd5)))};
  localparam signed [4:0] p10 = ((&(~(~^(~&(+((5'd30)<(4'd2)))))))<={4{(4'sd2)}});
  localparam signed [5:0] p11 = (2'd2);
  localparam [3:0] p12 = (-2'sd0);
  localparam [4:0] p13 = ((2'sd0)^~(-4'sd1));
  localparam [5:0] p14 = ((((~(4'd13))===(5'd15))<<{1{(-(&(3'sd1)))}})||{2{{1{(|(&(3'sd0)))}}}});
  localparam signed [3:0] p15 = {({(4'sd4),(3'sd2),(4'd1)}===((3'sd1)>(2'd1))),(5'd2 * {(4'd1),(5'd16),(2'd3)})};
  localparam signed [4:0] p16 = {2{(!(2'sd0))}};
  localparam signed [5:0] p17 = {3{(4'sd6)}};

  assign y0 = {(~|({p13,a0}-{p11,p11})),{(~&b2),(|p8),(b4&&p12)}};
  assign y1 = (((a1==a5)<=$unsigned(p4))&((b3<b1)%a3));
  assign y2 = (-(((a0^~p16)||(p12?b3:p11))?{2{{2{b4}}}}:{3{(p12<<p12)}}));
  assign y3 = (2'd2);
  assign y4 = ((~&((-3'sd0)!==(~^a2)))^~$signed((5'd1)));
  assign y5 = {3{(!p8)}};
  assign y6 = ((5'sd14)&&(-2'sd0));
  assign y7 = ((a1||a3)-(3'sd2));
  assign y8 = (2'd1);
  assign y9 = (|(~((p10?p15:p4)?(+p0):(^p9))));
  assign y10 = {(((p13<=p0)<={p5})<<$signed((+{b1,a5,p7}))),($signed({(~&p1),{p8,p3}})<=(+$unsigned({p3,p17,p10})))};
  assign y11 = ((a3===a3)>(a0>a5));
  assign y12 = (((|b1)!=$signed(b0))!==(^((^b4)<$unsigned(a5))));
  assign y13 = (5'd27);
  assign y14 = $signed({{(p16?p3:p3),{p16,p15},(p1?p11:p17)},({p3,p3}?{p2,p13,p6}:$signed((p12)))});
  assign y15 = (({3{(-p17)}}^~(~^((~|p11)||(-5'sd15))))-((2'd3)?{4{p9}}:(p17<=p14)));
  assign y16 = (((~^(-2'sd0))&&(&(5'd6)))>>>({b3,b0,a0}<<(5'd2 * (b2!==b1))));
  assign y17 = {{$unsigned(p4),$signed(b5)},{{2{a4}},{4{b3}},{2{p4}}}};
endmodule
