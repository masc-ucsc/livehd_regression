module expression_00219(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd3)?(5'sd0):(3'd7));
  localparam [4:0] p1 = ((6'd2 * (2'd2))?(|(5'd16)):((4'sd2)?(5'd9):(2'd3)));
  localparam [5:0] p2 = (5'd0);
  localparam signed [3:0] p3 = (~&(4'sd0));
  localparam signed [4:0] p4 = (((3'd2)?(-4'sd7):(-5'sd6))?((3'd4)>=(3'sd2)):((2'd2)|(-2'sd0)));
  localparam signed [5:0] p5 = {((4'd0)>(3'sd2))};
  localparam [3:0] p6 = {(~{(4'd4),(-2'sd1),(2'sd0)}),(~&{(5'd11)}),(&{(-2'sd1),(-4'sd0),(3'd7)})};
  localparam [4:0] p7 = (~(|(~|(~^(~(-(+(!(!(~|(&(&(~|(2'd3))))))))))))));
  localparam [5:0] p8 = ((-2'sd0)-(3'd5));
  localparam signed [3:0] p9 = ((3'sd1)>>>(~(((3'd2)<=(-4'sd4))||(|(4'sd4)))));
  localparam signed [4:0] p10 = {{4{((4'd12)>>(5'd14))}},({3{(3'd7)}}&&{2{(5'sd12)}})};
  localparam signed [5:0] p11 = ({(5'sd7)}<={(2'd0),(3'd5),(2'd0)});
  localparam [3:0] p12 = ((+((3'sd2)?(-3'sd0):(5'd22)))?((2'sd1)?(-3'sd0):(5'd20)):((3'd1)?(5'd6):(5'd7)));
  localparam [4:0] p13 = (((-3'sd0)>>(3'd1))>>((5'd10)^(2'd3)));
  localparam [5:0] p14 = ((4'd3)?(4'd15):(-5'sd0));
  localparam signed [3:0] p15 = ((~^((5'd23)|(4'd13)))||((5'd28)===(-3'sd0)));
  localparam signed [4:0] p16 = (3'd7);
  localparam signed [5:0] p17 = ((5'd2 * ((5'd31)?(2'd2):(3'd6)))<<<(((2'sd1)?(2'sd0):(4'sd7))<((5'sd2)?(-4'sd6):(4'd2))));

  assign y0 = ({p6,p11,b5}-(b1>=p14));
  assign y1 = (p11!=b3);
  assign y2 = ((|((a2==b1)>>(a5>>>a5)))+(~^((b3^p9)<=(a0>>a1))));
  assign y3 = (3'd5);
  assign y4 = ((~|(a1<=p8))>>>(p4!=p3));
  assign y5 = $unsigned(({2{p8}}));
  assign y6 = (&(!{1{{2{(&p10)}}}}));
  assign y7 = (&(4'd9));
  assign y8 = {2{{4{(a1|a3)}}}};
  assign y9 = (2'd1);
  assign y10 = ({(b3!=p12),(p13<<a1),(~p15)}?((p2?p16:p7)<={a0,a5,a1}):({p1,p4,p3}>(~p5)));
  assign y11 = (+(&((-(~^(((p15%p14)/p2)>>>((p14&&b2)<=(~&(^b2)))))))));
  assign y12 = ({1{{3{a1}}}}!=={1{(b3?a5:a2)}});
  assign y13 = (a2==p4);
  assign y14 = ((~&((~(b5==a0))>(p7+p4)))>>(~((p17&p9)-(p5>>>p17))));
  assign y15 = (({a5,b3}|(b4&&p1))<<{(-b0),{a0}});
  assign y16 = {({{2{b5}},(a0^b0),(b3===b2)}&({{{b3},{2{b5}}}}>>((a0?b4:b1)<<<(b3|b5))))};
  assign y17 = {3{(-2'sd0)}};
endmodule
