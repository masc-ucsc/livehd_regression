module expression_00494(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd4)/(-4'sd1));
  localparam [4:0] p1 = ({4{(2'd0)}}?{(-5'sd8),(2'd1),(5'sd7)}:((2'sd0)?(4'd14):(4'd6)));
  localparam [5:0] p2 = (~&(&(~^(~&(((4'd13)?(2'd0):(5'd16))?(+(5'd20)):{(2'sd0)})))));
  localparam signed [3:0] p3 = (~(2'd3));
  localparam signed [4:0] p4 = (&(-4'sd1));
  localparam signed [5:0] p5 = (-4'sd1);
  localparam [3:0] p6 = ({1{(3'd2)}}?{4{(2'd0)}}:(2'd0));
  localparam [4:0] p7 = ((((5'd14)!==(4'd13))+((2'd1)!==(-4'sd7)))+(+(+((2'sd1)%(-4'sd6)))));
  localparam [5:0] p8 = (~|(&(~({4{(2'sd1)}}===(4'sd2)))));
  localparam signed [3:0] p9 = (((-3'sd1)!=(5'sd14))?((-2'sd0)?(2'd3):(-3'sd0)):((-2'sd1)|(-4'sd1)));
  localparam signed [4:0] p10 = (6'd2 * ((5'd20)<=(5'd8)));
  localparam signed [5:0] p11 = {(3'd2),({(2'd3),(4'd10),(3'sd1)}>>(^(2'sd0)))};
  localparam [3:0] p12 = (&((5'd8)?(-2'sd0):(-4'sd2)));
  localparam [4:0] p13 = (|(~^(~&(|(^(~|(+(|(~(~(3'd5)))))))))));
  localparam [5:0] p14 = (+(~^(+(|{4{(&(-2'sd0))}}))));
  localparam signed [3:0] p15 = ((5'd11)<(5'd8));
  localparam signed [4:0] p16 = ((-3'sd0)+(-5'sd4));
  localparam signed [5:0] p17 = (&(((3'd1)==((4'd3)?(4'd5):(-5'sd7)))&(4'sd6)));

  assign y0 = ($signed((~^($unsigned($signed(b1))<<<(a0^~p4))))>>(($unsigned((4'd8))>>({4{p16}}>>>(p0>p8)))));
  assign y1 = ((|{1{(a3&b1)}})?((p6-p7)<(p3!=a1)):((a3)!=={1{b1}}));
  assign y2 = ($unsigned({1{{2{p6}}}})|(&(p5&p15)));
  assign y3 = ({a5,p15,a3}?(2'd0):(4'd7));
  assign y4 = ((~|$unsigned((|$unsigned(b2))))-(~^((~(b2>a0)))));
  assign y5 = {1{(((p14>>>p2)?{4{b5}}:(p2>=p11))?((+p11)<<<$unsigned(b3)):$unsigned({2{(p6)}}))}};
  assign y6 = (({2{p9}}||{4{a1}})?(5'd16):{1{((b0?p16:p5)<=(!b5))}});
  assign y7 = {3{({2{b3}}<<(a2===a4))}};
  assign y8 = (((p8?a0:p11)?(p12?p17:p0):(~&a3)));
  assign y9 = (~{(p1!=p16),{p14,b0},{p13,p16}});
  assign y10 = {(($signed((~|(~|b2)))^~(~^(b2||a0)))!=(^((~|((a0||b2)===(~^(&a2)))))))};
  assign y11 = (((p10<<p2)?(p16?b3:b0):(p10!=p0))||(^(~|((p5&p1)+(b5?p5:p9)))));
  assign y12 = {3{(b0>>>a1)}};
  assign y13 = {4{(-4'sd6)}};
  assign y14 = $signed($signed({3{(b3!==b5)}}));
  assign y15 = {((b3?p7:a4)?(b4>a1):(b4&b0))};
  assign y16 = ({3{a2}}>>>((p1?a3:p4)!=(p4?p7:p5)));
  assign y17 = $signed({{p2},{p14,b0},$signed(p10)});
endmodule
