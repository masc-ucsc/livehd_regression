module expression_00313(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((!(-5'sd12))^~((5'd10)<=(4'sd1)))^~(!(+{(-3'sd3),(4'd2),(3'd3)})));
  localparam [4:0] p1 = (4'sd4);
  localparam [5:0] p2 = ((3'd4)&(3'sd1));
  localparam signed [3:0] p3 = {3{{1{(((-5'sd13)==(-2'sd0))+(&(2'sd1)))}}}};
  localparam signed [4:0] p4 = (((-4'sd6)+(-5'sd12))&&((3'd0)==(5'd27)));
  localparam signed [5:0] p5 = (^(^((-2'sd1)==(3'd4))));
  localparam [3:0] p6 = ({3{(4'd14)}}>>((2'sd1)<=(2'd1)));
  localparam [4:0] p7 = ((4'd4)<(-2'sd1));
  localparam [5:0] p8 = (({(-3'sd0),(2'd1)}?(~(4'd3)):(~|(3'd0)))-{{((4'd2)!=(-3'sd1)),{(-5'sd3),(4'sd0),(-3'sd2)}}});
  localparam signed [3:0] p9 = ((-5'sd11)?(4'd4):(-3'sd3));
  localparam signed [4:0] p10 = (((3'd0)?(4'sd3):(-3'sd3))>>(&((5'sd12)||(3'd3))));
  localparam signed [5:0] p11 = (({(5'sd3),(-2'sd0)}||(&{(-4'sd1),(4'd8)}))>>{{4{(5'd0)}},((-5'sd13)<(2'd3))});
  localparam [3:0] p12 = {3{(((5'd11)&&(3'sd3))^~((5'd28)>=(5'd2)))}};
  localparam [4:0] p13 = (~(|(+(3'd7))));
  localparam [5:0] p14 = {4{((3'sd0)?(3'd0):(-3'sd2))}};
  localparam signed [3:0] p15 = ((3'd5)<<({1{((2'd1)&&(2'sd1))}}^(((3'sd1)>=(2'd0))===((4'd13)<=(-5'sd13)))));
  localparam signed [4:0] p16 = ((((2'sd1)&&(5'sd0))>=(~&{3{(5'd30)}}))&(~&({4{(2'd2)}}||((4'd15)<(-5'sd2)))));
  localparam signed [5:0] p17 = (|(3'd7));

  assign y0 = (!{p11,p10,p10});
  assign y1 = {3{{{a3,b0,b2}}}};
  assign y2 = (~|{3{((~p2)?(b1?a3:a0):(-5'sd9))}});
  assign y3 = (({b5})!=(~^(5'sd5)));
  assign y4 = (a5?b0:b2);
  assign y5 = (4'd2 * (!(&p13)));
  assign y6 = $signed(({1{(5'd22)}}));
  assign y7 = ((((~(~|b1))>((~a2)))!=(((!$unsigned(p17))^~(p12-p15)))));
  assign y8 = (b1>b1);
  assign y9 = (4'd4);
  assign y10 = ((((a4?a5:b4))?(~&$unsigned(b4)):$signed((b3?b3:b1)))===$unsigned(((b2?a5:a3)?(|(a1?b3:b3)):$unsigned((b0?b3:a2)))));
  assign y11 = (2'd3);
  assign y12 = ((b3?b2:b5)!==(b3-a5));
  assign y13 = {1{(~((4'd2 * (p6?p8:p2))<={2{(5'sd0)}}))}};
  assign y14 = (|(~^((b5!==a2)*((|p7)))));
  assign y15 = (-2'sd1);
  assign y16 = (!(!{(|(~&b3)),{a3,a1},{(^b5)}}));
  assign y17 = ({{a3,a3},(|p15),{a5}}>(-4'sd3));
endmodule
