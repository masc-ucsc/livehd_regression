module expression_00339(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd1);
  localparam [4:0] p1 = {1{(3'd1)}};
  localparam [5:0] p2 = (-(4'sd2));
  localparam signed [3:0] p3 = (((5'd2 * (4'd2))!==((-2'sd0)>>>(4'sd7)))+(((2'd0)<(2'd1))^{(3'd6),(-3'sd3),(-5'sd2)}));
  localparam signed [4:0] p4 = (((-5'sd5)?(-2'sd1):(5'd7))-(|(5'sd0)));
  localparam signed [5:0] p5 = (-(~(|(-3'sd2))));
  localparam [3:0] p6 = ((((2'd1)<<<(2'd1))<=(~^(~^(5'd16))))>>(((4'd7)^(2'sd1))<<((5'sd6)*(3'sd1))));
  localparam [4:0] p7 = ((-(|((2'd3)/(4'd10))))^(|(&(~|((4'sd6)^(4'd3))))));
  localparam [5:0] p8 = (~|(~|(~(~(2'sd0)))));
  localparam signed [3:0] p9 = (~^(-{4{(+((4'd1)?(2'd3):(-4'sd6)))}}));
  localparam signed [4:0] p10 = ((~&(5'd11))%(3'sd3));
  localparam signed [5:0] p11 = ((((-3'sd3)?(-2'sd1):(3'd2))>(~&(4'sd0)))?(~^(5'd2 * (2'd3))):((3'd5)?(4'd12):(2'd1)));
  localparam [3:0] p12 = (((4'sd1)|((2'd0)<<<(4'd10)))==(5'sd9));
  localparam [4:0] p13 = (((3'sd1)||(5'd13))?(~(5'd0)):(6'd2 * (2'd1)));
  localparam [5:0] p14 = ((~|{(5'd12),(2'sd0),(5'd27)})?{(&((3'sd1)>>>(2'd3)))}:{((2'sd0)?(4'd7):(4'd12))});
  localparam signed [3:0] p15 = (3'd7);
  localparam signed [4:0] p16 = ({3{((2'sd0)<<(3'sd2))}}|{1{({1{{4{(5'd13)}}}}>>>{{(4'd9),(2'd3)}})}});
  localparam signed [5:0] p17 = (-2'sd1);

  assign y0 = (2'd3);
  assign y1 = (2'd2);
  assign y2 = ({1{((p11&&p7)>>>(p5<<p1))}}<<<(&(~|(|((b3&b3)===(!a0))))));
  assign y3 = {1{$unsigned((&({a5,b1,b1}?((|p15)):$unsigned((a1?p0:b0)))))}};
  assign y4 = {({2{p16}}?{3{p8}}:(p6?p14:p11)),((p14?p3:p15)?(p1?p12:p6):(p15?p14:p0))};
  assign y5 = (b1|a2);
  assign y6 = ((b1>b5)?(a5&p11):(a1?p12:b3));
  assign y7 = (5'd2 * (2'd3));
  assign y8 = ((b3?p13:b4)?(p13?b0:a2):(p0?p15:p17));
  assign y9 = {1{((3'd5)?(~(~^$signed((5'sd4)))):((a1<=a5)||{1{{1{a4}}}}))}};
  assign y10 = (-3'sd1);
  assign y11 = {3{{1{b2}}}};
  assign y12 = (~&(4'sd7));
  assign y13 = {(~^{2{{1{(|b1)}}}}),{3{(~^$unsigned(a4))}}};
  assign y14 = (3'sd3);
  assign y15 = (b3);
  assign y16 = (5'd11);
  assign y17 = ({(&{p15,b5,b4}),(b1===b2),(^$signed(a2))});
endmodule
