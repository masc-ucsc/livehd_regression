module expression_00587(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd4)^~(((~(-3'sd2))!=(+(-3'sd3)))<<<(((2'd0)&(5'sd2))>>>(&(2'sd1)))));
  localparam [4:0] p1 = (5'sd6);
  localparam [5:0] p2 = (-4'sd3);
  localparam signed [3:0] p3 = (-(5'sd8));
  localparam signed [4:0] p4 = (~((2'd2)?(2'd0):(2'sd0)));
  localparam signed [5:0] p5 = (~|(~((|((4'd5)^(-4'sd1)))-((3'sd3)<<<(-4'sd1)))));
  localparam [3:0] p6 = (6'd2 * ((5'd25)+(2'd1)));
  localparam [4:0] p7 = (({(-5'sd2)}=={(3'd0),(3'sd0)})|(((2'd3)===(5'd15))<{(-3'sd0),(2'sd1)}));
  localparam [5:0] p8 = (|((^((5'd0)|(5'd16)))<<<((3'd1)?(3'd0):(-2'sd0))));
  localparam signed [3:0] p9 = ((+((2'sd0)!==(2'd3)))<{(^(-3'sd2)),{(2'd0),(3'sd0)}});
  localparam signed [4:0] p10 = {{{2{(4'sd5)}},(~^{(2'sd1),(4'sd3),(5'd25)})}};
  localparam signed [5:0] p11 = (3'd5);
  localparam [3:0] p12 = ({(4'd0)}^~((3'sd3)>>(3'd1)));
  localparam [4:0] p13 = (({4{(3'sd0)}}&{3{(5'd25)}})-({1{(4'd15)}}>>(~&(5'sd12))));
  localparam [5:0] p14 = (3'sd1);
  localparam signed [3:0] p15 = {((5'sd6)<(5'd23)),((4'sd3)<<<(-2'sd1))};
  localparam signed [4:0] p16 = {(&{{4{(-2'sd0)}},((5'd16)?(3'sd3):(5'd23)),((-2'sd1)?(-4'sd7):(-3'sd1))}),(-(^{(3'd0),(3'd4),(2'd3)}))};
  localparam signed [5:0] p17 = ((((-3'sd0)>=(-3'sd0))|((-3'sd0)===(4'sd7)))|({(-(-4'sd1))}<=((-2'sd0)^(5'sd14))));

  assign y0 = (+((^({p14,p14}^~{p10,p5,p13}))<<<({p8,p8,p7}&&{p8,p0,p3})));
  assign y1 = (((4'd14)|(b2?a4:p7))?{4{p12}}:{3{(~&a3)}});
  assign y2 = $unsigned(p9);
  assign y3 = (5'd8);
  assign y4 = (($signed((!b0))>>>(b1+p15))=={3{(~p17)}});
  assign y5 = (((-(b1-p13))>>>{(~&p16),(p1||p15)})^(((~&a4)!=(p12+p9))<(p17?a2:p12)));
  assign y6 = ((!((-4'sd6)|$signed(((a2==b0)===(b3|b4))))));
  assign y7 = {((a0+b1)<(a3>>p13)),(4'd6),((3'sd0)-{b0,b1,b4})};
  assign y8 = ((a4?a0:a5)===((b5?a0:a1)>(b2?b2:a2)));
  assign y9 = (-3'sd0);
  assign y10 = {((a0===b4)>>{b2,b2})};
  assign y11 = ((($unsigned((4'd14))==(p10<<<a4)))&&({(5'd2)}===(b5+a0)));
  assign y12 = ({p0,p6}!={p8});
  assign y13 = (5'sd4);
  assign y14 = (2'd3);
  assign y15 = (|(((-3'sd2)<(p3))>>>(4'd13)));
  assign y16 = ($unsigned((($signed(p11)-(p5^p0))>>>{1{{4{b0}}}}))>={1{{2{$unsigned((b2!==b4))}}}});
  assign y17 = ((~&((p10<<<p9)^~(a3!=p0)))^(~|(5'd16)));
endmodule
