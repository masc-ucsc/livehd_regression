module expression_00364(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(&(3'd7)));
  localparam [4:0] p1 = ((^(((3'd7)^(3'd6))<<((2'sd0)?(5'd17):(2'sd1))))>((+(4'sd3))?((-4'sd1)<<<(-5'sd2)):((4'd5)^(4'd6))));
  localparam [5:0] p2 = ({(5'd27),(3'sd0),(3'sd0)}+{((2'd2)|(2'd3)),((-5'sd15)?(-5'sd3):(2'sd1))});
  localparam signed [3:0] p3 = (-4'sd1);
  localparam signed [4:0] p4 = ((2'd2)?(-4'sd3):(-5'sd4));
  localparam signed [5:0] p5 = ((|{(5'd1),(-4'sd0)})^~(~&{(3'd0),(3'd1)}));
  localparam [3:0] p6 = (-{3{{(3'd3)}}});
  localparam [4:0] p7 = (~^((((-2'sd1)||(4'd15))<=(!(3'd3)))<((~&(2'd0))?((3'sd2)^(-2'sd1)):((2'd3)?(3'sd3):(3'd6)))));
  localparam [5:0] p8 = ((-2'sd1)?{(-3'sd3),(4'd1)}:{(3'd0),(2'd3)});
  localparam signed [3:0] p9 = (~(-2'sd1));
  localparam signed [4:0] p10 = (~&({(4'd0),(3'd4),(4'd1)}<=(&{(3'd7),(3'sd1)})));
  localparam signed [5:0] p11 = (~|(((2'sd1)>(4'd4))|((-5'sd13)^(-2'sd0))));
  localparam [3:0] p12 = (2'd3);
  localparam [4:0] p13 = (5'd15);
  localparam [5:0] p14 = ((|(2'sd1))<((4'sd4)<=(3'sd1)));
  localparam signed [3:0] p15 = (((5'd17)||(4'sd3))?((2'd2)!==(-4'sd2)):((-2'sd0)>=(-4'sd5)));
  localparam signed [4:0] p16 = (~|{3{(-{(-3'sd3),(-3'sd0)})}});
  localparam signed [5:0] p17 = (&((4'd2 * (2'd1))<<<{4{(4'sd4)}}));

  assign y0 = (^(~|((&p13)<<(a4+a2))));
  assign y1 = $unsigned(($signed(b3)==(a0?p17:b1)));
  assign y2 = {(3'd3),{4{p16}}};
  assign y3 = ({2{(b3===a4)}}<=(~&((a1?a4:p2)>>>{p10,a2,a4})));
  assign y4 = ({3{a3}}>>(|p9));
  assign y5 = (!((p14?p7:a1)?$unsigned((3'd3)):(p1>p16)));
  assign y6 = {{(b3?p8:b1),(a5&b5)},(5'd2 * (a2?p12:b1))};
  assign y7 = {2{(3'sd3)}};
  assign y8 = (((p11|p3)>>(p11<p0))||{(b2===b5),(p12+p11),{4{p1}}});
  assign y9 = $signed($unsigned($signed((4'd10))));
  assign y10 = ((p10)?(p17|p14):$signed(p17));
  assign y11 = $unsigned(($unsigned((($signed($signed($unsigned(((($unsigned($signed(p17)))))))))))));
  assign y12 = {4{{3{b0}}}};
  assign y13 = ((b0+b2)/a2);
  assign y14 = ($signed(p15)?(!p11):(-4'sd4));
  assign y15 = ($signed((3'd7))+{((b5<a0)^(b0<<<a2))});
  assign y16 = ({a2,a3}?(~a0):(~|b1));
  assign y17 = $signed({$signed({1{$signed({(&((p14<<<a3)|{p9,p8,a1}))})}}),((~|(!{p3}))|({a2,p11}+{3{b1}}))});
endmodule
