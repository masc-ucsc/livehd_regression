module expression_00314(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{3{(((4'd9)?(5'd20):(-4'sd4))>>>{1{(2'd0)}})}}};
  localparam [4:0] p1 = {2{(2'sd0)}};
  localparam [5:0] p2 = ((((5'd3)?(-5'sd8):(-5'sd0))>>>((-3'sd0)!==(2'd2)))&&({(5'd6)}>>>((3'd3)==(4'd7))));
  localparam signed [3:0] p3 = {{(-2'sd0),(3'd7),(5'd5)},((-5'sd7)>=(-2'sd1))};
  localparam signed [4:0] p4 = (4'd8);
  localparam signed [5:0] p5 = ((~((2'sd1)!==(5'sd11)))&&((5'sd10)&&(3'd5)));
  localparam [3:0] p6 = (4'd8);
  localparam [4:0] p7 = (((3'd7)/(4'd4))<=((5'd3)|(-2'sd0)));
  localparam [5:0] p8 = (~^(~|(4'sd1)));
  localparam signed [3:0] p9 = (+(-2'sd0));
  localparam signed [4:0] p10 = (((5'sd1)||(4'sd2))/(5'd2));
  localparam signed [5:0] p11 = ((((4'd15)>>(5'd27))<=((3'd5)>>>(3'd3)))|(^(((-4'sd1)&(5'd7))?((5'd2)!==(4'd10)):(+(4'd11)))));
  localparam [3:0] p12 = ((~((3'd6)?(2'sd1):(4'd6)))<{1{(~{2{(3'd5)}})}});
  localparam [4:0] p13 = ({2{((-3'sd0)!=(4'sd4))}}!==(-3'sd3));
  localparam [5:0] p14 = {(4'sd5),(3'sd1),(-3'sd0)};
  localparam signed [3:0] p15 = ((&(~|(~&(((3'd7)!=(4'd13))>>>(!(-2'sd1))))))<<(!((~|(~|(3'd2)))^(^(^(5'd28))))));
  localparam signed [4:0] p16 = (2'd2);
  localparam signed [5:0] p17 = (&(4'sd5));

  assign y0 = ((-3'sd0)>>(!(3'd4)));
  assign y1 = ((a2<=b2)||(a0?a0:b3));
  assign y2 = (+(~&({4{p10}}||(p3>>>b5))));
  assign y3 = {(&(|(^b3))),(^(a3===b4)),(~^(+(!b1)))};
  assign y4 = ({3{b0}}||({2{b3}}&&(3'd6)));
  assign y5 = (|(~$unsigned({(b1|p10)})));
  assign y6 = (&(((p3?p12:p5)?(4'd14):(p7!=p5))<<(5'd2 * (p12&p6))));
  assign y7 = (^((5'sd5)<<{p0,p10}));
  assign y8 = (b3!==b1);
  assign y9 = ({(!($unsigned(p10)>>>{p11,p6,p12})),(((^$unsigned(p6)))),{(p1<<<p16),(+p9),{p2}}});
  assign y10 = (~&{3{$unsigned($signed((p11?p4:p3)))}});
  assign y11 = $unsigned({(p1?p17:p0),(~^p14),(p6)});
  assign y12 = ((b0>a5)^(b4>>a5));
  assign y13 = (&($signed((a4>>>b3))<<<((4'd11)%p13)));
  assign y14 = ((-3'sd3)==={b5,b0,a2});
  assign y15 = ({2{((b1>>>p10)^~(p9?p11:a5))}}<<{1{($unsigned({3{a5}})?(a2<=p15):(p11?p2:b3))}});
  assign y16 = ((({4{a5}}===(b4!=b5))>>{4{p7}})||(4'd2 * {1{{1{p7}}}}));
  assign y17 = $signed((~|(&(~^$signed({{p13,a4,p16},{a5,p8},{p10}})))));
endmodule
