module expression_00960(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'sd3)!=(3'd1));
  localparam [4:0] p1 = (+(|(((-3'sd2)?(3'd0):(-2'sd0))?{(-4'sd1),(2'sd1),(5'sd5)}:((-2'sd1)?(2'sd1):(-3'sd0)))));
  localparam [5:0] p2 = ((~{(2'd2),(5'd28),(-3'sd0)})||(&(|((3'd0)?(5'd18):(3'd1)))));
  localparam signed [3:0] p3 = (&(^((((-3'sd3)-(5'sd12))%(5'sd15))^((^(3'sd3))||(6'd2 * (3'd3))))));
  localparam signed [4:0] p4 = {{(-2'sd0),(2'd2)}};
  localparam signed [5:0] p5 = {(((!((5'd14)^~(-4'sd5)))||(6'd2 * (2'd0)))=={{(3'd4),(4'd14),(2'd2)},((-3'sd0)>(5'd14)),(~&(-5'sd7))})};
  localparam [3:0] p6 = ((3'd3)?(2'd2):(5'd19));
  localparam [4:0] p7 = ((((3'd7)+(4'd3))%(3'd4))&&(((5'd5)!=(2'd0))>>>((5'd13)<<(3'd3))));
  localparam [5:0] p8 = (5'd2 * ((4'd1)===(3'd0)));
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = (-((^((+(3'd2))<<<((4'd4)!=(-4'sd7))))&{((2'd2)>>(-4'sd5)),(|(~&(2'sd0)))}));
  localparam signed [5:0] p11 = ((~|(^(-5'sd7)))==(2'd1));
  localparam [3:0] p12 = (|((~|(2'd1))?(~(4'sd0)):((4'sd4)?(4'sd0):(5'd12))));
  localparam [4:0] p13 = ((2'sd0)!=(2'd0));
  localparam [5:0] p14 = (-3'sd0);
  localparam signed [3:0] p15 = {{(5'sd11),(-3'sd2)}};
  localparam signed [4:0] p16 = ({1{(~^(~(4'sd4)))}}>=(|{3{(&(5'sd14))}}));
  localparam signed [5:0] p17 = {2{(4'sd7)}};

  assign y0 = (-({a3,b4}>>>(b5?p17:b5)));
  assign y1 = {({(~b0),(a1?b5:a3)}!==((~b1)?(a4>>>b1):(a2>a2))),(((+p15)?(a3===b2):{p5,p14,p11})^{3{(~p0)}})};
  assign y2 = ((((~b4)<=(~&b2))>=(~&{4{b5}}))>=(!(|(4'sd3))));
  assign y3 = ((-{2{(~^p12)}})^~({3{p16}}>>{4{p3}}));
  assign y4 = ((p3?p0:p2)<<(|(~&{2{p13}})));
  assign y5 = {4{((^(~|{4{p6}})))}};
  assign y6 = ($unsigned(p14)%p13);
  assign y7 = {{{b3,a2},{a4,a2}},{{{a1,a0}}},{p5,p12,b1}};
  assign y8 = {(-(~|(-{2{p8}}))),$signed({((4'd2 * a0)!=={2{a2}})}),({4{p12}})};
  assign y9 = {((b5?a0:b1)?{b3,p11,p9}:(-a2))};
  assign y10 = {2{((3'd2)?{4{p10}}:(2'd0))}};
  assign y11 = (((b3%p9)?(p8-p14):(p8*p13))>>((2'd1)||((b2%p13)<=(4'd0))));
  assign y12 = $unsigned((2'd1));
  assign y13 = ($unsigned((~&p17))<(a1!=a0));
  assign y14 = $unsigned($signed((^((~((p12==p15)))?(~&((~p15)<<$signed(p11))):(+(p6?p0:b5))))));
  assign y15 = {{{p4,p0},{p6,p17},{p13,b0,p7}},{{p13,p9},{a1,p14}}};
  assign y16 = (((b4+a3)+(a2===b2))!==((a0<=a5)===(&(b4!=b3))));
  assign y17 = (2'd3);
endmodule
