module expression_00661(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(4'sd2)}};
  localparam [4:0] p1 = (4'sd4);
  localparam [5:0] p2 = (~((~|((^(-2'sd1))|(^(2'sd1))))^~((~^(2'sd0))?(~(-5'sd1)):(!(2'd3)))));
  localparam signed [3:0] p3 = {1{(~|(^(~^{2{(-4'sd1)}})))}};
  localparam signed [4:0] p4 = {(((4'd12)>>>(-4'sd3))!=(^(4'd8)))};
  localparam signed [5:0] p5 = {(((|(4'd12))|((4'd14)>=(4'd6)))<<<(~^(|{((2'd0)!==(4'sd3)),((2'd2)||(4'sd5))})))};
  localparam [3:0] p6 = (|({(&(4'sd7)),((4'd10)<<(2'sd1)),((4'd13)===(-3'sd3))}>>(-(-3'sd0))));
  localparam [4:0] p7 = (-({1{(6'd2 * {1{((4'd10)<<<(4'd3))}})}}>>((4'sd6)<((-2'sd1)<<(-5'sd15)))));
  localparam [5:0] p8 = ((-2'sd0)?(5'd10):(4'd12));
  localparam signed [3:0] p9 = {{(5'sd14),(2'sd1)},{(-2'sd1),(3'sd1),(5'd3)}};
  localparam signed [4:0] p10 = ((5'sd4)^~(5'sd13));
  localparam signed [5:0] p11 = {3{{4{(-3'sd0)}}}};
  localparam [3:0] p12 = ((&(~((3'd4)?((2'd1)^~(4'sd0)):(^(5'sd6)))))===(^(~(6'd2 * (~|(~|(3'd7)))))));
  localparam [4:0] p13 = (|({3{(3'd0)}}>>>{2{(&(3'sd0))}}));
  localparam [5:0] p14 = (5'd5);
  localparam signed [3:0] p15 = (3'sd0);
  localparam signed [4:0] p16 = {{(|((4'd5)||(5'sd2))),{(|(3'sd1))}},(+(|{(2'sd1),(4'd5),(4'd8)}))};
  localparam signed [5:0] p17 = {3{{2{((-5'sd10)?(2'sd0):(3'sd2))}}}};

  assign y0 = ((~^(-5'sd9))^(5'd21));
  assign y1 = (~((-3'sd3)*(3'd2)));
  assign y2 = (~&(^((^(p12>=p3))/p2)));
  assign y3 = ({1{((~|(b0^a0))=={2{(p8<<b2)}})}}<<<{2{{4{a1}}}});
  assign y4 = (({b1,a0}!==(-2'sd0))?{2{(b1?p14:p15)}}:(~|(p1^a3)));
  assign y5 = (|$signed((-2'sd1)));
  assign y6 = ((b5?a5:a3)?((p3||b5)>=(b4!=a4)):((a3?p2:b5)>=(a0<=p9)));
  assign y7 = (3'd7);
  assign y8 = $unsigned(((5'sd8)==={(a3?a2:b5),{1{(b4?b4:b3)}},$signed((-3'sd0))}));
  assign y9 = (((a4||a4)!=$signed(b5))==={(-(b2-b1))});
  assign y10 = ({{(5'd2 * (p6|p1))}}-(((b1!==b5)|(p5>>p10))>>({p13,p7,p10}&{a3,p6})));
  assign y11 = ({1{((-{p14,p0,p12})&(p9^~p11))}}<={{3{(p14&p11)}}});
  assign y12 = (4'sd4);
  assign y13 = ((&(!(((a2-b0)<<(b2<=a3))>>((b5&&a1)===(-a3)))))===(^(4'd2 * (&(b2-b1)))));
  assign y14 = ({4{(|$signed(a4))}});
  assign y15 = {2{(4'd0)}};
  assign y16 = {1{{3{p5}}}};
  assign y17 = (((p9?p17:p14)||(p9>p16))-((p2?p1:p10)||(p15&&p11)));
endmodule
