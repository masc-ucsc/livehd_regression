module expression_00973(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'd1)?(2'd1):(3'sd3))?((-2'sd0)?(3'd6):(2'sd0)):(-5'sd2));
  localparam [4:0] p1 = ((|(4'sd4))||(~|((2'd0)|(3'sd3))));
  localparam [5:0] p2 = ((5'sd2)!=(4'sd0));
  localparam signed [3:0] p3 = {{((|(-3'sd1))?((3'sd3)?(4'd9):(2'd0)):((-5'sd12)?(5'd30):(5'd10)))}};
  localparam signed [4:0] p4 = (|((&(!(4'sd7)))||((4'd13)?(4'd5):(2'sd0))));
  localparam signed [5:0] p5 = (5'sd12);
  localparam [3:0] p6 = (&(~^(((3'sd3)?(4'sd5):(4'd14))>>(^(!((3'd4)?(-4'sd1):(-4'sd1)))))));
  localparam [4:0] p7 = (~^(&(~|(5'd6))));
  localparam [5:0] p8 = (|(|((^(~(-5'sd5)))^((-4'sd2)+(3'd4)))));
  localparam signed [3:0] p9 = (~&(~^(-(~^(-2'sd1)))));
  localparam signed [4:0] p10 = {1{(-4'sd0)}};
  localparam signed [5:0] p11 = (((2'sd1)?(3'd2):(4'd13))|(~^((2'd0)==(-4'sd5))));
  localparam [3:0] p12 = (5'd2 * {2{(5'd25)}});
  localparam [4:0] p13 = ((((2'sd0)>=(5'd8))>((3'd7)||(4'sd6)))||(((2'd1)<<<(3'd1))>((2'd0)<=(-2'sd0))));
  localparam [5:0] p14 = {((3'd1)?(2'd1):(-2'sd0)),{4{(5'd14)}}};
  localparam signed [3:0] p15 = ({(4'd4)}-(((3'd1)-(3'd1))&((5'd17)<(5'd20))));
  localparam signed [4:0] p16 = {3{((2'sd0)?(5'sd10):(5'd0))}};
  localparam signed [5:0] p17 = {{3{{(3'd2),(-2'sd0)}}}};

  assign y0 = (2'd1);
  assign y1 = (~^(+p15));
  assign y2 = (2'd2);
  assign y3 = (+(-(|(^((&{p17,a1,a3})<<<{(^{a2,p10})})))));
  assign y4 = (^(~&(-(5'd2 * {{a0,p6,a0}}))));
  assign y5 = (|(~(&(!{3{({4{a3}}?(a2?a1:a4):(~a5))}}))));
  assign y6 = (($unsigned(p5)==$unsigned(p0))&((6'd2 * b1)===(a4<<<b4)));
  assign y7 = {2{(~((!(a5>>a1))&(|(~^b0))))}};
  assign y8 = {2{((p11?p10:a1)|(b2^~p4))}};
  assign y9 = (&(3'sd2));
  assign y10 = ((((p1<p8)||(p9==p7))-((a0|a0)===(a1|a5)))>(((p4-p14)|(b4&&p2))==((a0>>>a0)!==(5'd2 * b0))));
  assign y11 = (2'd1);
  assign y12 = (-$unsigned((+$signed(b5))));
  assign y13 = ({3{p6}}?(a3?p3:b4):{a2,a3});
  assign y14 = (-4'sd4);
  assign y15 = (|(+({1{{2{(~&(2'd1))}}}})));
  assign y16 = (~|$signed((~(~|$signed((~^((!(3'd5))>>>(|$unsigned((a4|p2))))))))));
  assign y17 = (a2?a3:a2);
endmodule
