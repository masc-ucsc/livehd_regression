module expression_00546(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(^{(4'sd3)}),(((-4'sd5)?(2'sd0):(4'd8))?(2'sd0):((3'd2)?(4'sd5):(5'd31)))};
  localparam [4:0] p1 = ((((5'd30)^(2'd1))>>>((4'd14)>>>(4'd15)))!==(((3'd6)<<<(2'd3))?((-2'sd0)>>>(-4'sd4)):((3'd5)!=(5'd21))));
  localparam [5:0] p2 = (~{2{{3{{(-5'sd14),(3'd3)}}}}});
  localparam signed [3:0] p3 = (-2'sd1);
  localparam signed [4:0] p4 = ({(2'd2),(5'd2),(-3'sd0)}<<<{4{(-5'sd10)}});
  localparam signed [5:0] p5 = (((4'd2)?(2'd2):(4'sd2))?((5'd21)?(2'd1):(2'd1)):((-4'sd5)?(-2'sd0):(4'sd4)));
  localparam [3:0] p6 = {3{(~|(-3'sd3))}};
  localparam [4:0] p7 = ((|(!(~|(-5'sd10))))&&{{4{(4'd5)}},{1{(2'd2)}}});
  localparam [5:0] p8 = ((|((-3'sd3)^~(3'd7)))?((-4'sd6)^~(-3'sd1)):((5'd5)*(4'sd5)));
  localparam signed [3:0] p9 = ((^(~^((-3'sd1)<((3'd3)>>>(4'd6)))))<<(-2'sd0));
  localparam signed [4:0] p10 = ((~^(+{(2'd2),(-4'sd3),(-4'sd3)}))!=(~|((5'sd7)?(-2'sd0):(-3'sd2))));
  localparam signed [5:0] p11 = ({3{(4'd6)}}?{1{((3'd3)?(5'd2):(-5'sd15))}}:(|(&((2'sd1)?(5'sd7):(3'd3)))));
  localparam [3:0] p12 = (2'd1);
  localparam [4:0] p13 = ({{(5'd11),(-2'sd0)},{((5'd23)>>(3'sd3))}}^~(((4'sd0)^~(5'd22))|{3{(5'd23)}}));
  localparam [5:0] p14 = {((-2'sd1)>(4'd13)),((-4'sd5)|(3'd7)),{(5'sd13),(-5'sd11)}};
  localparam signed [3:0] p15 = {3{(4'd12)}};
  localparam signed [4:0] p16 = (-3'sd2);
  localparam signed [5:0] p17 = (+((((-4'sd5)!==(-5'sd6))/(-3'sd0))^(~|((-3'sd1)!==(5'sd10)))));

  assign y0 = ((-(5'd2 * (~^(a0&a1))))===(((b1)^(^a1))&($signed(b3)?(b2):(a0?b3:a3))));
  assign y1 = ($unsigned({(((a3<a5)>{(b5==a5)}))})==={{b1,b2},{$signed(a3)},(b0-b1)});
  assign y2 = (((b3>=b1)>>>(a1!==a2))&&(!(a5|a3)));
  assign y3 = (-((^{(~|{$unsigned(p7),$unsigned(p15)}),(~&(~|$unsigned({p12}))),$unsigned((|(-{p13,p0})))})));
  assign y4 = ((~((p17>>>a4)?(&a4):(a0^~a0)))&&((b0?a4:a3)|(b5?p9:b5)));
  assign y5 = (((5'd3)?(~^a0):(p5^a2))?((+a0)?(p13&p17):{4{a3}}):{1{{4{p6}}}});
  assign y6 = (!((4'sd6)==(4'sd5)));
  assign y7 = (-2'sd0);
  assign y8 = (~{(|(+(&(!a4)))),(|({b2}<<(|a4)))});
  assign y9 = ((b5<p14)?(5'd27):(p12?a3:a3));
  assign y10 = (^(~^a2));
  assign y11 = {4{(^{p6,p12,p9})}};
  assign y12 = (~(5'd4));
  assign y13 = {3{((a3>>>a4)>>{3{b3}})}};
  assign y14 = (p8==p3);
  assign y15 = $unsigned((~|(~|$unsigned(((~(^(+{b1,b3,b0})))<(-$signed((!(^a5)))))))));
  assign y16 = {4{b3}};
  assign y17 = {2{(+{1{((b3+p13)&{1{(&b2)}})}})}};
endmodule
