module expression_00380(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-2'sd1)?(4'sd5):(2'd1))&&((-3'sd1)*(3'd3)))&&((|(3'sd1))?(+(3'd0)):(~&(4'sd7))));
  localparam [4:0] p1 = (((~^((4'sd2)?(5'sd12):(-2'sd1)))<<(~((4'd15)?(2'd1):(4'sd4))))>>>(!((+(~(4'd13)))*(~|((2'd1)?(-5'sd2):(2'sd1))))));
  localparam [5:0] p2 = {(~((-3'sd3)-(4'sd3))),(&((2'd3)<<(5'd15))),{(3'd2),(5'd10),(5'd15)}};
  localparam signed [3:0] p3 = (~&(4'd12));
  localparam signed [4:0] p4 = ((((-4'sd2)|(2'd0))>((5'd25)!==(4'd1)))?(|{(^(-4'sd6))}):{{(2'd3),(-3'sd1),(-3'sd3)}});
  localparam signed [5:0] p5 = (4'd2 * ((2'd0)>(5'd1)));
  localparam [3:0] p6 = (((3'd3)&&(-3'sd1))?((4'd14)%(4'sd3)):((3'd6)>=(-4'sd2)));
  localparam [4:0] p7 = (((-4'sd5)-(2'd1))<<(4'd2 * (4'd13)));
  localparam [5:0] p8 = ((~|{3{(-3'sd0)}})?(((5'sd3)!==(-5'sd8))>((4'sd6)?(5'd4):(-4'sd0))):{3{((5'sd3)>>(3'd7))}});
  localparam signed [3:0] p9 = (((-((5'd10)==(3'sd0)))<<<{(-2'sd0),(4'sd5),(-5'sd3)})>>(~(5'd2)));
  localparam signed [4:0] p10 = (-5'sd9);
  localparam signed [5:0] p11 = ({((3'd0)&(5'd20)),{2{(-4'sd2)}}}?(((-5'sd7)&(-3'sd3))=={4{(2'sd0)}}):{3{{2{(4'd4)}}}});
  localparam [3:0] p12 = ((&((4'd4)?(3'sd1):(4'sd4)))?((-5'sd10)!=(-5'sd3)):(5'd9));
  localparam [4:0] p13 = ((~|(3'sd2))^~(&(4'd11)));
  localparam [5:0] p14 = (3'd3);
  localparam signed [3:0] p15 = ((5'd30)*(3'd6));
  localparam signed [4:0] p16 = {((~^(5'd28))?((-5'sd6)<(2'd0)):((-2'sd1)==(-2'sd1)))};
  localparam signed [5:0] p17 = ((4'd10)^(3'd0));

  assign y0 = {4{(b2?b0:a2)}};
  assign y1 = ((!((b3?a4:p6)!=(-3'sd2)))?(~|(~^(b2?b1:p4))):((+p8)?(!b2):(|b0)));
  assign y2 = ((($unsigned(b2)<<<(-2'sd0))>=(-3'sd0)));
  assign y3 = ({{4{{b4}}}}==={{2{a5}},{4{b4}},{(a0>=b3)}});
  assign y4 = (3'd0);
  assign y5 = (4'd8);
  assign y6 = (|p12);
  assign y7 = {(~^(((p5?p9:b4)==($unsigned($unsigned(p2))))&&(!(|((b2?a0:a2)?(a5&&b1):(b2>>>b0))))))};
  assign y8 = (((-5'sd7)?(5'd2 * b2):(b2?a1:a2))===((a0===b5)?{1{a3}}:(b4-a1)));
  assign y9 = ({3{p3}}!={p17,p10,p9});
  assign y10 = $signed({2{(((p5?p5:p5)&&((a5===a3))))}});
  assign y11 = ({(3'd0),(b2==p2),(|b4)}||((^(3'd5))>=(p3>=p0)));
  assign y12 = (^((p0<<<p2)!=(b2===b0)));
  assign y13 = ($unsigned((4'sd4))>>$unsigned(((&(~&p13))|(b1?b0:a0))));
  assign y14 = ((4'd5)+(a4<<a2));
  assign y15 = (((&(^(p11)))&&((b3|p9))));
  assign y16 = {3{{2{(5'd2 * a0)}}}};
  assign y17 = (&(!(4'd2 * (^(5'd20)))));
endmodule
