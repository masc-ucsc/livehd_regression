module expression_00051(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(5'd0)}};
  localparam [4:0] p1 = ((((3'd3)?(-4'sd2):(3'd2))*(3'd3))?((^(3'd1))?((5'd28)!=(4'd12)):((4'd8)>>>(5'd20))):(5'd10));
  localparam [5:0] p2 = ((3'd0)|(2'd0));
  localparam signed [3:0] p3 = {{2{(3'd2)}},{(2'sd1),(2'd1)},{(5'sd13),(3'd5)}};
  localparam signed [4:0] p4 = ((3'd2)-(4'sd3));
  localparam signed [5:0] p5 = (!((~&(~^((~^(4'sd1))>(-3'sd2))))>((~^(-3'sd2))?(2'sd1):((5'sd13)<<(2'd3)))));
  localparam [3:0] p6 = ((((5'sd15)!=(2'd1))==((2'sd1)&&(5'd16)))>=(2'd1));
  localparam [4:0] p7 = ((3'd2)>(5'd27));
  localparam [5:0] p8 = {2{(~|{4{(5'sd10)}})}};
  localparam signed [3:0] p9 = (|(~&((2'd1)&&(-4'sd2))));
  localparam signed [4:0] p10 = ((2'd0)?(5'd13):(-5'sd10));
  localparam signed [5:0] p11 = (3'd4);
  localparam [3:0] p12 = (~&(~&(~&(|(+(~&(~^(+(~^(-4'sd1))))))))));
  localparam [4:0] p13 = (^(!{(~&(5'sd11))}));
  localparam [5:0] p14 = ((((2'sd1)<=(5'd30))>(~&(4'd5)))-{((3'd3)<<(-2'sd0)),{(3'd3),(2'sd0)}});
  localparam signed [3:0] p15 = {4{(3'd7)}};
  localparam signed [4:0] p16 = ((-3'sd0)&(((-3'sd0)!==(2'd1))?((-5'sd10)&&(2'd1)):(6'd2 * (3'd4))));
  localparam signed [5:0] p17 = {3{((5'sd5)<(4'sd5))}};

  assign y0 = (((b5&b3)>=(b3%a1))&((a4<<<a1)||(b3/b2)));
  assign y1 = (~&{1{a2}});
  assign y2 = {(p15-a0),(p15?p9:p5),{p10}};
  assign y3 = (~(~(&(&{p4,p5}))));
  assign y4 = (|(^({(-p11),{3{p6}},{a3,p3}}?(-(a1?p2:p4)):($signed(p6)?{4{p5}}:{a4,p14,p17}))));
  assign y5 = ((^(~^{{2{b0}},{2{p17}}}))|(~{(~^p12),(-4'sd2)}));
  assign y6 = (&(~^(~&(-(!$signed($signed((b5|a5))))))));
  assign y7 = (2'd0);
  assign y8 = (|(~$signed((-{2{((b4?a4:a1)?(a1&a1):(a0>=p8))}}))));
  assign y9 = (b2|p3);
  assign y10 = (-2'sd1);
  assign y11 = (&(!(~^((~|(~|(|(!b3))))|(~((4'd2 * a2)===(2'sd1)))))));
  assign y12 = $unsigned(($signed((p17?p14:p7))?((p14?p16:p6)?(p7||p15):(b3?p12:p6)):((p14*p8)?(p15):(p6?p17:p4))));
  assign y13 = ((^(~|(((p2?a2:p13)!=(!b3))+((b1?p11:p2)*(&p9)))))>>((~&((p3>>a3)<<<$signed(a1)))!=((p17==p15)<=(&p4))));
  assign y14 = ({2{(-2'sd0)}}<<{3{{3{a2}}}});
  assign y15 = ((a4^b4)?(-5'sd12):(a3?p3:b5));
  assign y16 = (({1{{4{b3}}}}<<<(a2>a4))^~((p14?a0:p13)?(a0>>b1):(p15-p12)));
  assign y17 = (~^(~&(!($unsigned((^(~(~|($unsigned((-(!(~(2'd1))))))))))))));
endmodule
