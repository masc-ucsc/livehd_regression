module expression_00006(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&{1{((((4'sd7)-(2'd0))&&(~^(5'd4)))==((-5'sd11)?(4'd1):(-3'sd1)))}});
  localparam [4:0] p1 = (3'd1);
  localparam [5:0] p2 = (({(5'd3),(4'd4)}+{(5'sd6)})!==(|(|(~^(4'd4)))));
  localparam signed [3:0] p3 = (~^(|(5'sd0)));
  localparam signed [4:0] p4 = ((((5'd30)<<<(-5'sd0))?((4'sd4)?(-3'sd1):(5'sd3)):(&(-5'sd11)))?((4'd2 * (3'd7))?{1{(5'd20)}}:((4'd13)^(5'd6))):(^(((2'd3)?(-4'sd0):(4'sd5))<<((-2'sd0)>(3'd0)))));
  localparam signed [5:0] p5 = (-(2'd3));
  localparam [3:0] p6 = ((5'd18)<(((5'sd11)^(3'd2))>(-3'sd2)));
  localparam [4:0] p7 = (4'd2 * (3'd1));
  localparam [5:0] p8 = (~&{4{{4{(-3'sd1)}}}});
  localparam signed [3:0] p9 = ({2{(4'd1)}}<=(3'sd1));
  localparam signed [4:0] p10 = (~|(^((~^(-5'sd7))+(~|(-4'sd3)))));
  localparam signed [5:0] p11 = (3'sd3);
  localparam [3:0] p12 = ((-2'sd1)===(5'd3));
  localparam [4:0] p13 = (2'd0);
  localparam [5:0] p14 = (((5'sd4)/(3'd0))%(-4'sd2));
  localparam signed [3:0] p15 = ((~({2{(2'd3)}}?((-4'sd4)-(-2'sd0)):(6'd2 * (2'd2))))<<<{3{(4'sd0)}});
  localparam signed [4:0] p16 = (-3'sd0);
  localparam signed [5:0] p17 = {(4'sd2),(4'sd7),(-4'sd4)};

  assign y0 = (a5!==a0);
  assign y1 = (({3{p0}}&{2{a1}})<<{1{(~&{p15,p1,b4})}});
  assign y2 = {({a1,p2,a1}^~(+(a5?b5:p9)))};
  assign y3 = ((~|($signed({b4})^~(p14?b1:p6)))?{$unsigned($signed((a2?p5:b1)))}:((p11?p9:a0)?(b5?p1:b1):(b2)));
  assign y4 = (((~&a4)!=={3{a0}})+{4{a5}});
  assign y5 = $unsigned(((a2?p9:p12)));
  assign y6 = $signed((-3'sd0));
  assign y7 = ((-((^a2)<=(b2<=p0)))&{3{{3{p14}}}});
  assign y8 = {{(5'sd8),{4{b4}},(p4?b5:a5)},((!b1)?(a5?a1:a3):(a5?b4:p11)),{{3{b0}},(4'sd4),{b3}}};
  assign y9 = {4{{p14,p14,a3}}};
  assign y10 = (5'd24);
  assign y11 = (5'd20);
  assign y12 = $signed({(((-4'sd4))?{p9,a4}:(5'sd9)),(((~|(p0&&b1)))|{(p12?b3:p0),(p17?p12:b1)})});
  assign y13 = (((p13?p10:p10)&&({p0}>=(p8^p15)))<(~&(3'd3)));
  assign y14 = ((~^(~|(~^p6)))&((p5!=p12)^~(!p14)));
  assign y15 = (^$unsigned((($signed(p9)?(p9?b1:b4):(a1?b3:p8))?((&(!{p13,a3,b4}))):(+(-{p13,p13,a2})))));
  assign y16 = ((p16&&p14)?(p8):(&b5));
  assign y17 = (p0?p12:b5);
endmodule
