module expression_00848(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{1{((4'd1)?(4'd7):(4'd9))}}}};
  localparam [4:0] p1 = ((~^(+(|(2'd3))))===((~|(2'sd0))+(+(2'd1))));
  localparam [5:0] p2 = (|(3'sd2));
  localparam signed [3:0] p3 = ({(-2'sd0),(5'd21),(-3'sd3)}?({(-4'sd2)}^((4'd14)?(3'sd2):(2'sd1))):((-5'sd0)^~((-4'sd4)?(4'd9):(-4'sd1))));
  localparam signed [4:0] p4 = (((3'sd2)===(4'd12))<<<((3'sd2)===(3'd0)));
  localparam signed [5:0] p5 = {(({(4'd3),(-3'sd2)}>>(^(5'd5)))<((-(5'd16))==((5'sd1)===(-2'sd0))))};
  localparam [3:0] p6 = {3{(4'd9)}};
  localparam [4:0] p7 = {{((4'd11)<<<(3'd1)),((-5'sd14)>=(4'd9)),(~^(~&(5'd27)))},(((2'd0)^(-2'sd0))?(&((4'd3)<<(4'sd1))):(^((5'sd7)?(-4'sd0):(4'sd2))))};
  localparam [5:0] p8 = (5'd5);
  localparam signed [3:0] p9 = {({(5'd25),(-2'sd1),(2'd2)}==={(5'sd15),(3'd1),(5'd7)})};
  localparam signed [4:0] p10 = ((&(5'sd14))?{2{(-4'sd5)}}:((3'd5)>=(5'd6)));
  localparam signed [5:0] p11 = ((^{{(-3'sd0)},((-5'sd14)?(2'sd0):(4'd9))})+{({(5'd29),(2'sd1)}||{(2'd0),(4'sd3)})});
  localparam [3:0] p12 = ((4'd2)<=(5'd2));
  localparam [4:0] p13 = (~&{4{{(-5'sd9),(4'd0),(4'd3)}}});
  localparam [5:0] p14 = ((((5'd31)<<<(-4'sd6))||((-3'sd2)|(3'sd0)))+{3{{1{(5'd9)}}}});
  localparam signed [3:0] p15 = (((~|(5'sd14))!==(&(3'd1)))?(((5'd21)?(5'd19):(2'sd0))-((5'sd4)!==(5'd7))):(5'd2 * ((3'd1)^(2'd0))));
  localparam signed [4:0] p16 = {4{(+(-3'sd3))}};
  localparam signed [5:0] p17 = (((3'd7)^~(-3'sd0))!=={3{(-3'sd2)}});

  assign y0 = ({{{(^(b0!=a3))},((-b1)>>{1{b2}})}}||{3{(b5?a4:a0)}});
  assign y1 = ((-2'sd1)<=((-4'sd7)||(a0^~a4)));
  assign y2 = ($unsigned((5'd6))==(&(~|(+(2'd3)))));
  assign y3 = {1{{2{{3{p4}}}}}};
  assign y4 = ((a3?b5:p2)<<(a1?p8:p6));
  assign y5 = (-5'sd4);
  assign y6 = ((((5'd18)|(~|p0))||(!{b4,p14}))+((p16?p8:p2)?(b1<=a1):(p12^b1)));
  assign y7 = (|(((&(~b3))+({4{p16}}))+(~|(3'd0))));
  assign y8 = {4{(-$signed($signed(p17)))}};
  assign y9 = {3{b1}};
  assign y10 = ($unsigned({2{(p8)}})!=(|($unsigned(a1)>>(a3===a0))));
  assign y11 = (((p17-p6)<=(p16?b3:p13))?((p11?a1:a5)>>(~^p11)):((&p13)*(^p4)));
  assign y12 = (+({(2'd3)}<<<((a4?b5:a0)>(3'd1))));
  assign y13 = (((+b1)==={2{b2}})&&{3{p12}});
  assign y14 = (-(~^(^(-((~|$signed((^a1))))))));
  assign y15 = ((5'sd9)?(3'd2):((-5'sd11)>=(p15||a0)));
  assign y16 = (+(~|b2));
  assign y17 = ((((b0<<p10)<<$unsigned((b3===b5)))==((b5-p5)<(a0^~p1))));
endmodule
