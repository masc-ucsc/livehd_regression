module expression_00554(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((-(3'sd2))%(-4'sd4))>>(~&((4'sd0)>>>(2'd3))))+(((2'd1)^(-4'sd2))?((2'd1)*(2'd3)):((2'sd0)&(3'sd3))));
  localparam [4:0] p1 = ((-(~^(3'sd2)))<<<((-4'sd0)+(5'd22)));
  localparam [5:0] p2 = ({((-5'sd6)!==(4'sd1)),(^(5'sd14))}|(-3'sd3));
  localparam signed [3:0] p3 = (3'sd1);
  localparam signed [4:0] p4 = (((!(4'd15))?(-(-3'sd3)):(&(2'd3)))?(~&(~^(!(+(4'd9))))):((~^(5'd4))-(+(-3'sd0))));
  localparam signed [5:0] p5 = ({2{((3'd2)?(2'd3):(-2'sd1))}}>>>(|{2{{1{(-3'sd1)}}}}));
  localparam [3:0] p6 = (({1{(-5'sd10)}}>{3{(5'sd5)}})>>>{{(5'd8)},((5'd23)<=(4'd5))});
  localparam [4:0] p7 = (((3'sd1)?(-5'sd12):(3'd2))?((2'sd1)?(3'd4):(2'sd1)):((-2'sd1)/(-2'sd0)));
  localparam [5:0] p8 = ((~(^{(3'd6),(-4'sd2),(3'sd1)}))!=(-(~|{(~(2'sd1))})));
  localparam signed [3:0] p9 = {((3'd2)+(-3'sd2))};
  localparam signed [4:0] p10 = (!((((4'sd6)<<(3'd4))>(^((5'd22)==(2'd0))))<=((&(~^(2'd3)))!=(+((2'd3)^~(5'd29))))));
  localparam signed [5:0] p11 = ((~(-((5'sd3)>=(-2'sd1))))<<<({(2'd2),(5'd20)}<<(6'd2 * (4'd12))));
  localparam [3:0] p12 = ({(3'd7),(2'sd0),(5'sd5)}>>>(!(+(~^(-5'sd12)))));
  localparam [4:0] p13 = ((-2'sd0)==(5'd7));
  localparam [5:0] p14 = ((4'd14)<<(2'sd0));
  localparam signed [3:0] p15 = {3{(~&(~&((4'd12)>=(3'd5))))}};
  localparam signed [4:0] p16 = (~(((4'd0)+(5'sd3))>((3'sd2)?(4'd6):(-2'sd1))));
  localparam signed [5:0] p17 = ((((3'sd0)==(3'd0))>>((-4'sd4)|(4'sd7)))===((&(3'd1))-((3'd1)&&(2'd0))));

  assign y0 = (~&(!(-(a3?p8:b3))));
  assign y1 = (&(({(p0-p12)}^(^(p15<=p5)))?((-(p12&p5))&&$signed((p16?p2:p0))):((p12<p4)||($unsigned(p6)))));
  assign y2 = (((b0&a2)==={2{a0}})&({1{{3{b0}}}}>>>(p8^p10)));
  assign y3 = (~^{(&(-(b4>p3)))});
  assign y4 = ((~((p10<p13)?(b5&a5):(+b2)))<<<((b1^~b4)!==(a0<<<b0)));
  assign y5 = (5'd14);
  assign y6 = ({(p15||p16),(6'd2 * b2),(p1^p0)}<<((p4!=p4)>>{p0,p10,p3}));
  assign y7 = ((2'sd0)<{2{p0}});
  assign y8 = {3{(b5?p7:b4)}};
  assign y9 = ($unsigned(((a1>=b2)+{b2,b4,b2}))!=$unsigned(($unsigned({a3,b3,a4}))));
  assign y10 = (((6'd2 * p7)&&(p7|p2))&$signed((p12?p12:p15)));
  assign y11 = ((5'd31)/a2);
  assign y12 = {((~|(3'd7))?(~&{p1}):(~|{4{p1}})),(!((~p13)?(|b5):{1{b1}}))};
  assign y13 = (!(&((|a5)?{1{p12}}:{1{b2}})));
  assign y14 = {(&((~^b0)?(a1<=p9):{b4,a0,b1})),((a5?b4:a4)>(~^(+b3)))};
  assign y15 = ({2{((a5&&p16)<<(|b5))}}|({3{a4}}<((-p13)<(b5!==a3))));
  assign y16 = (&{{(a2!==b2),(a0>>p12)},((p1!=p17)?(p6?a1:a1):{3{a4}}),{2{(b0|b0)}}});
  assign y17 = ((2'd3)?(-(4'd11)):(p14^~p13));
endmodule
