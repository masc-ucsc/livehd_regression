module expression_00290(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{{(4'd5),(5'sd2),(-4'sd7)},((5'd30)?(5'sd1):(-2'sd1))},(((3'sd3)?(5'd11):(3'd4))<<<((3'd3)?(3'd6):(3'd7)))};
  localparam [4:0] p1 = (-3'sd3);
  localparam [5:0] p2 = (+((5'sd14)^~((-5'sd0)!=((3'd6)?(-5'sd5):(2'd1)))));
  localparam signed [3:0] p3 = {{((5'd7)+(3'd0)),((4'd13)+(-4'sd4))},(-{(-(3'd0)),{(4'sd5),(3'd6),(2'd1)}}),{(!(5'd4)),(!(-3'sd2)),((2'sd0)||(-4'sd4))}};
  localparam signed [4:0] p4 = (~&{3{(-(4'd9))}});
  localparam signed [5:0] p5 = ((^(-(-(2'd1))))^(2'd3));
  localparam [3:0] p6 = ((6'd2 * ((4'd2)<(4'd7)))<(((4'sd1)<<(5'sd8))>>>((-2'sd1)<<(4'sd1))));
  localparam [4:0] p7 = (!(~|(|(~|((2'd2)<(-2'sd1))))));
  localparam [5:0] p8 = (4'd15);
  localparam signed [3:0] p9 = {2{(3'd4)}};
  localparam signed [4:0] p10 = ((6'd2 * (4'd11))>>((2'sd1)||(4'd14)));
  localparam signed [5:0] p11 = (6'd2 * {(4'd12),(3'd4),(3'd0)});
  localparam [3:0] p12 = (~{3{(((3'd1)!=(5'sd8))||(4'sd0))}});
  localparam [4:0] p13 = ((-5'sd12)?(5'sd13):((5'd2)?(5'd28):((5'sd0)?(3'd7):(-2'sd0))));
  localparam [5:0] p14 = {3{(4'sd1)}};
  localparam signed [3:0] p15 = ({(4'sd1),(4'd10),(3'd0)}?((4'd2)?(2'd3):(2'sd0)):{{(3'd4),(3'd7),(3'sd3)}});
  localparam signed [4:0] p16 = ((((5'd18)?(3'sd2):(-5'sd5))&&(5'sd3))<=((-3'sd1)?(4'd10):(2'd2)));
  localparam signed [5:0] p17 = (((~(5'd30))||((4'sd4)?(3'd5):(-3'sd0)))?(~^((-3'sd0)?(3'd0):(4'd15))):((~(3'sd0))?(-(-4'sd1)):((2'sd1)&&(3'd7))));

  assign y0 = (|$signed($unsigned(((~(3'sd2))!=$unsigned($unsigned((~p10)))))));
  assign y1 = (3'd4);
  assign y2 = (|(4'd8));
  assign y3 = {1{(&(((|b2)&&(a1!=b2))!==(!((a2|a2)&&(-a0)))))}};
  assign y4 = ((~{1{((4'd12)^(5'd4))}})>=(5'sd10));
  assign y5 = (~|(p12^~p11));
  assign y6 = (!((|(~&$unsigned((~^b5))))>>>((~|p6)?(b5|p12):(p7>>>p14))));
  assign y7 = ((~&{1{{b5,p3,p7}}})^~{4{a1}});
  assign y8 = $signed(((!(p4>=p16))%a4));
  assign y9 = (4'd1);
  assign y10 = {2{((&{4{p2}})<{3{p3}})}};
  assign y11 = {2{(3'sd2)}};
  assign y12 = (5'd14);
  assign y13 = (({b4,p2}>(p9&&a4))>>>{(-p1),(+p11),(p0?a1:p1)});
  assign y14 = $signed((&$signed(((p15)/b0))));
  assign y15 = (4'd8);
  assign y16 = {(b4!==b4),{4{p14}}};
  assign y17 = ({{{p14}},(p17?p9:p6),(b2?p15:a3)}^~((p12<<<b1)?(b3!=a0):(!(|p15))));
endmodule
