module expression_00584(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd1);
  localparam [4:0] p1 = (({3{(5'd11)}}&&((-3'sd2)&(-5'sd5)))<<{4{((-3'sd0)>>(2'd3))}});
  localparam [5:0] p2 = (|(4'd10));
  localparam signed [3:0] p3 = (~&(~&{{(-5'sd12),(4'sd6)}}));
  localparam signed [4:0] p4 = {(((4'd6)===(-4'sd6))+{(3'sd3)})};
  localparam signed [5:0] p5 = (({1{(-5'sd11)}}?{(3'sd3),(3'd4)}:((3'd2)?(5'd28):(4'sd0)))!==({(4'sd2)}?{(2'd1),(5'd21),(3'sd3)}:{(-4'sd3),(4'sd0)}));
  localparam [3:0] p6 = {4{((-2'sd1)?(-4'sd4):(4'd2))}};
  localparam [4:0] p7 = (2'sd0);
  localparam [5:0] p8 = (~|(2'd0));
  localparam signed [3:0] p9 = (-(-3'sd3));
  localparam signed [4:0] p10 = {1{{2{(3'd2)}}}};
  localparam signed [5:0] p11 = (~^((-(2'd3))?((-5'sd11)^~(4'sd5)):(~&(3'd0))));
  localparam [3:0] p12 = ((4'd1)?(5'sd9):(5'd26));
  localparam [4:0] p13 = {3{((2'sd0)<<<(2'd1))}};
  localparam [5:0] p14 = ((~^((4'sd4)>>>(3'sd3)))^(((2'sd1)<(2'sd1))>>>(-(4'sd1))));
  localparam signed [3:0] p15 = ({(4'd14),(|{4{(4'sd1)}})}<=(6'd2 * {((5'd31)<<(4'd10))}));
  localparam signed [4:0] p16 = {1{(-(~|(|(!({3{(5'sd7)}}?(-5'sd12):{2{{4{(-3'sd3)}}}})))))}};
  localparam signed [5:0] p17 = (-{((4'd8)<<(5'sd2)),{(-2'sd0),(2'd1)}});

  assign y0 = (((~^(a3?p15:b0))&(-3'sd1))?(4'd2 * (5'd21)):((^(~b1))^(2'd3)));
  assign y1 = {{{1{({2{p16}}+(p8!=p10))}}},{{p0},(p16==p10),{p4,p0,p0}},({4{p9}}!=(p17|a2))};
  assign y2 = ({($unsigned(p15)>=(-5'sd9)),$signed({$unsigned(a0),{a0}})}^($unsigned({{b4,b2},(4'sd6)})===$signed($unsigned($unsigned((b5+b5))))));
  assign y3 = (a0===a0);
  assign y4 = ((4'd2)<=(((4'd2 * p7)-(b4?p1:b3))==$signed(((a5>>p6)))));
  assign y5 = {3{(p3&&p6)}};
  assign y6 = (-4'sd2);
  assign y7 = (-4'sd3);
  assign y8 = ((a2&&a0)?(a1?a1:b3):(-4'sd0));
  assign y9 = {({p7,b5,a1}<<<{4{a2}}),(!(^(a4^a5)))};
  assign y10 = (((4'd2 * p12)=={a3})<<((^p1)<=(|a3)));
  assign y11 = ((4'd13)^~(4'd10));
  assign y12 = (|(!((~(&(b5?a5:a2)))?(&(b4/b5)):(a3?a3:a2))));
  assign y13 = (~&(&(5'd30)));
  assign y14 = (p3?b2:p0);
  assign y15 = (^{4{{3{(b3-a3)}}}});
  assign y16 = ({{1{{4{a5}}}}}^~{(+(~&a5)),{2{b0}}});
  assign y17 = (-2'sd0);
endmodule
