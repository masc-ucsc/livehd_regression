module expression_00552(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(!((5'd9)?(3'sd3):(2'd0)))}};
  localparam [4:0] p1 = (({(4'd12),(5'd15)}==={{(-5'sd15),(2'd1)}})-(((3'd5)?(5'sd9):(5'd7))-((-2'sd0)>=(5'sd7))));
  localparam [5:0] p2 = {3{((~(4'd8))?((4'sd3)>>(2'd0)):{(5'sd15),(5'd29)})}};
  localparam signed [3:0] p3 = ({4{(2'd0)}}<=((2'sd1)||(4'sd2)));
  localparam signed [4:0] p4 = (((|(3'd2))<((5'sd7)||(5'sd13)))!=((!(-5'sd5))+(^(-3'sd1))));
  localparam signed [5:0] p5 = ((4'd8)>=(5'd22));
  localparam [3:0] p6 = (2'sd1);
  localparam [4:0] p7 = ((5'd6)<(2'd0));
  localparam [5:0] p8 = {{4{((3'sd1)===(2'd0))}}};
  localparam signed [3:0] p9 = {(!((3'sd0)>>(3'd0))),{1{((4'sd1)>(4'd2))}},{1{(~(2'd3))}}};
  localparam signed [4:0] p10 = (-(~&(4'd15)));
  localparam signed [5:0] p11 = (&(5'd14));
  localparam [3:0] p12 = (3'sd1);
  localparam [4:0] p13 = (((4'sd3)>((4'd1)?(-3'sd3):(-5'sd6)))<<(6'd2 * (2'd3)));
  localparam [5:0] p14 = ((((2'd2)>(4'd11))>=((5'd14)&(2'sd1)))<<<{{(4'd9),(3'sd3)},((4'd11)!=(2'd1))});
  localparam signed [3:0] p15 = (~(3'sd2));
  localparam signed [4:0] p16 = ((~(-(((5'd24)&(3'sd0))-(|(4'd3)))))!=(~{(-(-3'sd2)),((3'd1)<=(3'd1)),((3'd5)!=(4'd10))}));
  localparam signed [5:0] p17 = ((2'sd0)>=(-4'sd0));

  assign y0 = (($unsigned(b0)<{a4})>>>((b0?b5:p2)>>>$unsigned(a0)));
  assign y1 = (!p17);
  assign y2 = {3{((b4>>a4)!==(b0^~a4))}};
  assign y3 = $signed($signed({{3{a0}},(b1),{b4}}));
  assign y4 = (-(^(&({a2}^(!a4)))));
  assign y5 = {2{{2{(p14^p0)}}}};
  assign y6 = (4'sd7);
  assign y7 = {{3{{a3}}},(4'd2 * {p0,b2,a1})};
  assign y8 = $unsigned($unsigned((|(+$signed((^(~&p16)))))));
  assign y9 = (4'd1);
  assign y10 = $signed((((-b3)?(5'sd2):$unsigned(p7))?((-2'sd0)+(p14?p15:b4)):(|((p13<=a1)+$unsigned(p6)))));
  assign y11 = {3{{2{(|a1)}}}};
  assign y12 = (&(((!($unsigned(p8)!=(b3&p3))))^~((a4|a1)!=(&(~|a4)))));
  assign y13 = (p7^~b1);
  assign y14 = ({(~&(a1>>>b1)),{b1,a5}}?({{a2,a3}}<<<(2'd1)):{(~a3),(~^a5),(b2|a0)});
  assign y15 = {{2{($unsigned({p4})<<(p3&a1))}}};
  assign y16 = (^{4{(~^b3)}});
  assign y17 = ((3'd3)-(3'd3));
endmodule
