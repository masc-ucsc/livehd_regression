module expression_00531(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd0)>>{(&(4'd0))})!=(4'd3));
  localparam [4:0] p1 = (^({(2'd2),(2'sd0),(5'sd9)}?((2'd0)?(-2'sd1):(-2'sd0)):(~(~(2'd3)))));
  localparam [5:0] p2 = ((5'd0)?(-4'sd3):(-4'sd7));
  localparam signed [3:0] p3 = (({(4'd4)}^~(^(4'd2)))||(|(|((-5'sd11)?(2'd3):(5'd17)))));
  localparam signed [4:0] p4 = {(~|(|{(~(~{(2'sd0),(5'sd0),(3'd4)})),{(~{(-3'sd0)})}}))};
  localparam signed [5:0] p5 = (~^(-((^(!(4'd12)))?(!((3'd1)?(2'd3):(2'sd0))):((5'sd10)?(-5'sd4):(4'd13)))));
  localparam [3:0] p6 = ((((4'd3)-(5'sd12))+(&(5'd14)))>>>{{1{(-4'sd1)}},(&(4'd13))});
  localparam [4:0] p7 = ((4'd4)?(-3'sd1):(^(-5'sd12)));
  localparam [5:0] p8 = (((+(-2'sd0))?((4'd5)?(3'sd0):(2'd2)):(&(-5'sd6)))!=(((3'd7)?(-2'sd0):(2'sd1))>>>((-4'sd4)?(2'd2):(3'd0))));
  localparam signed [3:0] p9 = (&(((3'd4)!=(3'd6))>((4'd10)>>>(3'd2))));
  localparam signed [4:0] p10 = ((((3'sd0)&(-2'sd1))!=((2'sd0)?(2'd1):(2'd2)))?(((2'sd1)<<<(5'd4))?{4{(4'sd4)}}:((-3'sd0)|(5'd13))):(^{2{((2'd1)!=(-3'sd1))}}));
  localparam signed [5:0] p11 = (&((-5'sd9)<(3'sd1)));
  localparam [3:0] p12 = {({4{(-5'sd5)}}?(^(2'sd1)):((4'sd1)&&(5'd17))),(|{((2'd3)==(3'd3)),((3'd4)?(2'sd1):(5'd8))})};
  localparam [4:0] p13 = ({1{((5'd22)&&(-5'sd13))}}!={1{((-2'sd0)<=(4'd0))}});
  localparam [5:0] p14 = ({(&((3'd0)>(4'd8)))}>>(!(2'sd0)));
  localparam signed [3:0] p15 = (^(+(~|(^(-(^(!(+(|(~|(|(-(~|(~|(~&(5'sd5))))))))))))))));
  localparam signed [4:0] p16 = (((4'd13)!=(-(2'd1)))-(&((|((2'sd1)*(-4'sd0)))>=((3'd4)||(-2'sd1)))));
  localparam signed [5:0] p17 = {{(5'd2 * (3'd0)),{(-5'sd2),(2'sd0),(4'd3)},(~(-2'sd0))},{2{(~^((4'd15)==(-4'sd0)))}}};

  assign y0 = {1{({4{{1{b2}}}}>>{(~(p5!=b5)),{(p4>p8)},{1{(~p1)}}})}};
  assign y1 = (((a1&p6)>>>(p7<<<p8))&((2'sd0)>>>(2'sd1)));
  assign y2 = (4'd9);
  assign y3 = (4'sd4);
  assign y4 = ({(~&(p12?p16:p9)),(a2?b3:a2),$unsigned((p10+p8))}==($unsigned($signed(p16))?(5'd12):(-5'sd10)));
  assign y5 = ((((^p15)&(a0>>>p12))>=((a3>>>p15)!=(^p2)))<<(((a5>>b3)&(a0^~p3))||((a4<p9)<=(p15>a5))));
  assign y6 = $signed(((!((|b1)==(5'd2 * b2)))?((!b4)&(p5?a1:b5)):((3'd7))));
  assign y7 = ((~(5'd24))^((!(a0===b2))<(5'sd15)));
  assign y8 = {2{(+$signed((~&(~&({4{a5}}<<{3{p4}})))))}};
  assign y9 = (3'd7);
  assign y10 = (3'sd3);
  assign y11 = (b3?a2:p1);
  assign y12 = (((b3<<<a4)<=(a0<b3))&(4'd2 * {b1,b0}));
  assign y13 = (5'd2 * (4'd14));
  assign y14 = (($unsigned({{b5}})));
  assign y15 = ((!{((~&p16)^(~b4)),(p15?p12:p4)})==((((a5!==a5)===(b0==a0)))!==($signed((a1?b4:b3)))));
  assign y16 = (p15&p0);
  assign y17 = (((p15?a5:b5)?(b5?a3:p0):{2{b1}})?((~|p13)?(b2?a2:p14):(-a3)):(-(a2?b5:p0)));
endmodule
