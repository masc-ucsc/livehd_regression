module expression_00471(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'sd1)||(3'd3))>>((5'sd8)/(2'd1)))?(((-4'sd3)>>(-5'sd15))+((4'd2)?(2'd0):(-5'sd10))):(((4'sd4)<=(3'd7))||((5'sd8)?(2'd3):(2'd0))));
  localparam [4:0] p1 = ((-(5'd6))<=(~^(5'd25)));
  localparam [5:0] p2 = {{2{{(-4'sd2),(-4'sd4),(2'd3)}}},{1{(((5'sd13)==(5'd4))^~(+(3'd2)))}}};
  localparam signed [3:0] p3 = ((((5'd30)^(-3'sd3))&((3'd3)?(2'd1):(2'sd0)))===(((2'sd0)-(-5'sd12))&&(!((2'sd0)>=(2'd2)))));
  localparam signed [4:0] p4 = ((^((3'sd1)<(3'sd2)))?((2'd1)?(5'sd15):(2'sd0)):((-3'sd2)!=(3'd7)));
  localparam signed [5:0] p5 = (((-3'sd3)?(-4'sd7):(4'd7))?(|((-5'sd8)?(5'd19):(5'd3))):(~&((5'sd12)?(2'sd1):(3'd1))));
  localparam [3:0] p6 = ({1{(4'd11)}}<<<((-2'sd1)<<(5'd18)));
  localparam [4:0] p7 = (({2{(5'sd9)}}?((4'd1)>=(-2'sd0)):(&(3'd5)))?{1{((-3'sd0)?(5'd19):(3'sd1))}}:((~(2'd3))?((-4'sd1)?(3'd4):(-4'sd1)):((2'sd0)&(2'd0))));
  localparam [5:0] p8 = (3'd3);
  localparam signed [3:0] p9 = {{((5'sd6)?{(5'd1),(5'd13)}:(5'd28))},(3'd4)};
  localparam signed [4:0] p10 = ((((5'd16)&(2'd0))>((5'sd5)!==(-4'sd5)))^(((2'd1)<<<(5'd31))===((-4'sd3)>=(-2'sd0))));
  localparam signed [5:0] p11 = {(4'd0),(4'd14),(-3'sd3)};
  localparam [3:0] p12 = ({(-4'sd3),(2'd2),(-4'sd5)}?(-{4{(2'sd1)}}):{(5'd7),(-2'sd0)});
  localparam [4:0] p13 = {4{((3'd7)>(-2'sd1))}};
  localparam [5:0] p14 = ((((4'd1)?(4'd14):(-3'sd3))>=(5'd11))>=({(3'sd3),(2'd1)}>>>((3'd5)<=(4'd6))));
  localparam signed [3:0] p15 = (5'd18);
  localparam signed [4:0] p16 = (3'sd1);
  localparam signed [5:0] p17 = (((|(4'd2))>(|(3'd4)))-((-5'sd12)<=((3'd0)%(3'd2))));

  assign y0 = {4{(~^((p6>>p0)!=(-p11)))}};
  assign y1 = (((p3?p14:p17)?(-(p15+p4)):(p6?b1:a1))>((~|(p12?b2:b4))?(~^(a2<=p2)):(p12-a3)));
  assign y2 = (((!a4)&&(b3?b1:b2))!=={((~&b5)>>>(+a4))});
  assign y3 = ((~(^b4))|(p7==b1));
  assign y4 = (3'd0);
  assign y5 = ((4'd0));
  assign y6 = (~^(&(~^(-5'sd1))));
  assign y7 = {(5'd2 * (5'd1)),(-2'sd1)};
  assign y8 = {{p3,p16},$signed(p0)};
  assign y9 = (+a4);
  assign y10 = {4{{a3,a0}}};
  assign y11 = (~&(((-(~&{4{b5}}))>((!a4)===(-b2)))^{2{(~&{4{p6}})}}));
  assign y12 = {({p0}!=(p13?p6:p13)),((p17?p11:p13)?(b1+p17):(p3<=p3)),{(~^(|{p0,p16,p2}))}};
  assign y13 = ((^{1{(-{(a1|p16),{4{b3}}})}})-({4{p16}}||((~|p3)?{4{p0}}:(p7!=p11))));
  assign y14 = (!$signed({2{b2}}));
  assign y15 = (~({4{(a3?p13:p0)}}));
  assign y16 = {{a5,p16},(p9>=a5),(b4-p9)};
  assign y17 = ((|(a3!==a5))===(~|(+(a1*a2))));
endmodule
