module expression_00594(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd3);
  localparam [4:0] p1 = (6'd2 * (4'd2 * (2'd1)));
  localparam [5:0] p2 = (6'd2 * ((3'd5)+(4'd3)));
  localparam signed [3:0] p3 = (~|(5'd22));
  localparam signed [4:0] p4 = (-5'sd10);
  localparam signed [5:0] p5 = ((3'sd2)>>{1{(-(4'd7))}});
  localparam [3:0] p6 = {{(~^(|{3{((3'd5)!=(3'sd0))}}))}};
  localparam [4:0] p7 = ({2{((2'd2)>(4'd8))}}<<<(-((4'd4)>=(3'sd3))));
  localparam [5:0] p8 = (~(!(~(5'd2))));
  localparam signed [3:0] p9 = (((-2'sd0)?(5'sd4):(5'sd2))?(2'd2):(2'd0));
  localparam signed [4:0] p10 = (~&(-(+(|(+(~(|(~^(^(-(+(!(&(|(-2'sd1)))))))))))))));
  localparam signed [5:0] p11 = (|(2'd0));
  localparam [3:0] p12 = ((^(3'd1))?(!((-2'sd1)?(4'd14):(-3'sd1))):(-2'sd1));
  localparam [4:0] p13 = {1{{2{({3{(2'd0)}}!==(|(+(5'sd12))))}}}};
  localparam [5:0] p14 = (|(~|(4'd2 * ((5'd9)%(5'd7)))));
  localparam signed [3:0] p15 = (((~^(-5'sd15))?((5'd1)>>>(4'd6)):((4'd7)>(4'd7)))?(((3'd0)^(3'sd1))%(3'sd0)):(((4'd13)>>>(4'd7))|((5'd19)>(5'sd2))));
  localparam signed [4:0] p16 = {4{{1{{4{(4'd14)}}}}}};
  localparam signed [5:0] p17 = (3'd0);

  assign y0 = (-{({p14}?{b2,p9}:(|a3)),((&a5)?{a3,p0,b4}:(~^p16)),(~^(~&{(p14?b2:a0),(-p14)}))});
  assign y1 = $unsigned(((~(2'd2))===({4{b0}}!==(-3'sd2))));
  assign y2 = $signed($signed(((b3<a2)?(~(p12?b1:b1)):((|p17)))));
  assign y3 = (&(~&(((|a4)?(a4?a1:a2):(-b3))-({3{p3}}-(b3?b0:b2)))));
  assign y4 = (((p8?p12:p10)?(p7>p15):(p14?p17:p6))<=((p4<p10)?(p2^a1):(b4?p5:p8)));
  assign y5 = ((b4?a5:b3)<<<(~&(b4?b3:a1)));
  assign y6 = ({2{b2}}+{4{a2}});
  assign y7 = {1{{1{{((p15<=p6)>={2{p10}}),{4{(a2<<<p13)}},{3{{p11,p8,b4}}}}}}}};
  assign y8 = (((~&(~^a0))?(a4&b1):(b2<<b2))!==(((b1?b3:b4)!==(!b1))^(b5?b5:a0)));
  assign y9 = ((4'sd3)&((p9^~p8)>{1{b5}}));
  assign y10 = (-3'sd2);
  assign y11 = (4'd2);
  assign y12 = (((~(!(&p6)))<<(~(p0|p13)))<<(((&b0)<<<(~|b0))===(|(b1!==b3))));
  assign y13 = ((2'sd0)?(-4'sd3):{1{a0}});
  assign y14 = ({({{a4,b1,a2}}>(4'd8))}<$signed((4'sd5)));
  assign y15 = $unsigned($signed((-5'sd15)));
  assign y16 = {3{(a4!=a2)}};
  assign y17 = ((~&((a5!==a0)===(5'd18)))<=($signed($unsigned(b1))&(a5===a4)));
endmodule
