module expression_00070(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(&{{(^(2'd2)),(~&(5'd13)),(-(-2'sd0))},{(+(4'sd3)),{(2'd2)}},(+{(~(4'd6)),((4'd14)&(-4'sd1))})}));
  localparam [4:0] p1 = ((((2'd2)?(2'd1):(2'd2))>(5'sd12))?(2'sd0):((4'd13)?(5'sd11):(4'd11)));
  localparam [5:0] p2 = (|(~&(~(~|(+(3'd6))))));
  localparam signed [3:0] p3 = (2'd1);
  localparam signed [4:0] p4 = (-5'sd12);
  localparam signed [5:0] p5 = (-(+(&(^((4'd2 * (5'd19))<<(~^((5'd17)!=(3'sd1))))))));
  localparam [3:0] p6 = (~^(((-3'sd3)<<(3'd4))^(~&(~|(5'd3)))));
  localparam [4:0] p7 = {(5'sd11)};
  localparam [5:0] p8 = (((-2'sd1)-(-3'sd2))!==(({(5'd20)}>(2'd3))&&(((2'd3)^~(2'd3))<=((4'sd0)^~(-2'sd0)))));
  localparam signed [3:0] p9 = (|(~^(~&(+(~|(+((!(5'sd2))!=((-5'sd10)^~(-3'sd0)))))))));
  localparam signed [4:0] p10 = ((3'sd3)^~(~&(2'sd0)));
  localparam signed [5:0] p11 = (((4'd14)|(2'd3))/(2'sd1));
  localparam [3:0] p12 = {4{(3'd3)}};
  localparam [4:0] p13 = (+((3'd7)||({(-5'sd5),(5'd17)}^~((3'd4)<=(2'd0)))));
  localparam [5:0] p14 = (((-2'sd1)?(-4'sd4):(3'd6))&&((4'd6)?(4'd5):(3'd0)));
  localparam signed [3:0] p15 = ((((3'd3)^(3'd2))>>((5'd31)+(5'sd1)))+({(5'd20),(-5'sd3),(4'd0)}-((5'sd6)?(3'd0):(4'sd5))));
  localparam signed [4:0] p16 = ((&((4'sd4)-(5'd30)))/(-3'sd1));
  localparam signed [5:0] p17 = (-4'sd2);

  assign y0 = (!(5'd23));
  assign y1 = {{2{{(!p11),(p12<<<p5),(p16<<<p3)}}}};
  assign y2 = (5'd2 * a0);
  assign y3 = ((p3%p6)^~(-2'sd1));
  assign y4 = (((p17<<p17)*(3'sd2))>>((4'sd1)*(-2'sd0)));
  assign y5 = ((2'd2)?({3{b0}}^(b5^a5)):(5'd12));
  assign y6 = ((3'd6)/b1);
  assign y7 = (|((p0<<p12)*(5'd16)));
  assign y8 = ({3{p7}}^~(p17||b5));
  assign y9 = ((3'sd3)>=$signed((5'd2)));
  assign y10 = ({3{$signed({1{$signed({2{a0}})}})}});
  assign y11 = (~({(p1&p10),(!p8),{3{p15}}}||(~|{2{{2{p3}}}})));
  assign y12 = (~&a1);
  assign y13 = (~|(((a2||b0)<(-a5))>>>{1{({2{b3}}^~(b5>>p1))}}));
  assign y14 = ((3'd7)&(~^((3'd7)^(b0===a1))));
  assign y15 = ((~|$unsigned(($signed(((a1*b5)<<(+(a5>>>b5)))))))^$signed((((b5&&a4)/a0)<<<((5'd2 * a0)))));
  assign y16 = {a2,a0};
  assign y17 = {1{{2{p2}}}};
endmodule
