module expression_00950(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~{(~|(|(~|{{2{(&(4'd10))}}})))});
  localparam [4:0] p1 = (-(-5'sd11));
  localparam [5:0] p2 = {((5'd16)?(2'sd1):(3'd3))};
  localparam signed [3:0] p3 = (!(({(2'd1),(4'sd1),(2'sd1)}^~{(4'd11),(4'd1),(3'sd1)})||(2'sd0)));
  localparam signed [4:0] p4 = (&(|(-3'sd0)));
  localparam signed [5:0] p5 = (!(~|(-3'sd2)));
  localparam [3:0] p6 = {4{((5'd22)?(-5'sd10):(-4'sd3))}};
  localparam [4:0] p7 = ({((5'd4)===(5'd29)),(~|((5'd29)==(-3'sd3)))}>>>((-(~(5'sd2)))||(-4'sd4)));
  localparam [5:0] p8 = (~|{1{(+(|({(~(2'sd1)),{(-4'sd6),(-5'sd0)}}!=(!(~{(-3'sd3)})))))}});
  localparam signed [3:0] p9 = (+(~&((2'd3)<=(3'd6))));
  localparam signed [4:0] p10 = {2{(((4'sd7)|(3'd1))-((2'sd0)>>(2'sd0)))}};
  localparam signed [5:0] p11 = {((~(5'd8))^((2'd1)>(4'd10))),{(((-3'sd0)>>>(2'd2))|{(-2'sd0),(5'sd3),(5'd4)})},(^{1{(~^{(4'd4),(2'sd0),(5'd16)})}})};
  localparam [3:0] p12 = ((~|((!(2'sd1))?(!(5'sd11)):(~&(3'd4))))||((|(&(4'd14)))==((5'sd12)*(-2'sd0))));
  localparam [4:0] p13 = {3{(5'd16)}};
  localparam [5:0] p14 = {2{((-2'sd0)&(2'sd0))}};
  localparam signed [3:0] p15 = (3'd0);
  localparam signed [4:0] p16 = ((4'd11)?(^(((3'd2)!==(5'd8))>>>(5'd7))):(((5'd18)+(3'sd2))?((4'd9)>>>(3'd6)):(~|(5'd23))));
  localparam signed [5:0] p17 = (2'd0);

  assign y0 = ({({b0,a4,a3}>>(b2!==a0)),({b0}<={b5})}<<((b0-b0)?(b0==a0):{(b1?a5:a2)}));
  assign y1 = {3{((|b3)|(a1))}};
  assign y2 = ({2{a5}}===(~^b1));
  assign y3 = (2'd1);
  assign y4 = {4{(3'sd2)}};
  assign y5 = ({{((p7>>a4)>>>(a1-p7))}}==(!(~&(^{{b4,p11},(!(~|a3))}))));
  assign y6 = (4'd2 * (p1?b2:a2));
  assign y7 = (b2<<p17);
  assign y8 = ((p2/p14)^$unsigned(b4));
  assign y9 = $signed(((a2?p12:p10)&(p5==p15)));
  assign y10 = {1{({$unsigned(p16)}?({3{p3}}):$unsigned($unsigned(p10)))}};
  assign y11 = (((b3===a1)&(4'd10))!=((a5<=b3)<=(~^b2)));
  assign y12 = (&{4{a1}});
  assign y13 = ({4{(^p17)}}<<((p7^~p11)>>((~&p10))));
  assign y14 = {2{p6}};
  assign y15 = (((p11+p0)^~$unsigned(p4))<<{4{p10}});
  assign y16 = (-(!({(4'sd7)}^(3'sd1))));
  assign y17 = ({1{{1{(4'd3)}}}}-(^(3'sd1)));
endmodule
