module expression_00191(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-5'sd0);
  localparam [4:0] p1 = (&(((+(-4'sd6))>(~(4'd9)))>=(~^(-3'sd1))));
  localparam [5:0] p2 = ({1{(5'd2 * ((4'd9)?(4'd6):(5'd13)))}}?({2{(4'sd1)}}!==(|(4'sd6))):((~|(5'd19))?((2'sd1)|(2'd2)):((2'd2)<=(3'sd0))));
  localparam signed [3:0] p3 = ((((5'd4)&(2'd0))&((2'd3)<=(5'd22)))-(((4'sd1)|(-2'sd1))<((5'd4)===(-3'sd3))));
  localparam signed [4:0] p4 = {2{{4{(5'd3)}}}};
  localparam signed [5:0] p5 = (~|(~&(3'sd2)));
  localparam [3:0] p6 = {(!(|{(-3'sd2),(-3'sd0)})),(~|(~^((4'd9)<<(3'sd1))))};
  localparam [4:0] p7 = {(5'd28),((~&(-4'sd6))>>(!(5'd22))),(3'sd3)};
  localparam [5:0] p8 = (~(({(4'sd4),(2'd1)}>((2'sd0)&&(5'd19)))!==((~|{(-5'sd3),(-3'sd3)})&&(3'sd0))));
  localparam signed [3:0] p9 = (3'sd0);
  localparam signed [4:0] p10 = (+(-(!(-(|{2{(!{4{(3'd3)}})}})))));
  localparam signed [5:0] p11 = ((5'd5)<=((-5'sd13)?(-5'sd5):(3'd2)));
  localparam [3:0] p12 = ((^(&((2'sd0)?(2'd0):(5'd13))))|(!(((-4'sd2)<<(3'sd2))<(-(2'd2)))));
  localparam [4:0] p13 = (!{4{(-3'sd3)}});
  localparam [5:0] p14 = ((~|((-4'sd7)<=(3'd0)))%(5'd30));
  localparam signed [3:0] p15 = {1{{2{{4{(4'sd4)}}}}}};
  localparam signed [4:0] p16 = (((2'd2)?(5'd1):(-4'sd6))?(-5'sd3):(4'd14));
  localparam signed [5:0] p17 = {{(-2'sd0),(3'd4),(5'd28)},((3'd1)>>>(-3'sd3)),{(|(-5'sd12))}};

  assign y0 = (((5'd7)?{(+b5)}:(-3'sd3))=={(-4'sd1),{(~&(b2?b0:a5))}});
  assign y1 = (((p12<=p3)?{4{p17}}:{4{p0}})^((-2'sd0)|(p5?p13:a5)));
  assign y2 = (~((~|(5'd2 * (b1?p6:p0)))^~((4'd0)||(-(b5?b2:a4)))));
  assign y3 = (((p4?b0:a3))^$unsigned($signed(a1)));
  assign y4 = ((3'd7)!=(-4'sd7));
  assign y5 = ({4{a0}}^~{{1{p17}},{a4,a0}});
  assign y6 = (|(~^{{{(|p0)},{a3,b1},{b4,a2,p12}}}));
  assign y7 = (5'sd10);
  assign y8 = ($signed(((a0?p1:a3)-$unsigned(a3)))?((p8?p17:p6)?(p10?p4:p14):(a4?p5:b4)):((p12>>>p12)?(p6==p3):$unsigned(p3)));
  assign y9 = $unsigned($signed(($signed(($unsigned((($signed($signed($signed($unsigned($signed(($unsigned(b2)))))))))))))));
  assign y10 = {(((b4>=b1)>=(~(b4?b1:b3)))?((3'd4)+(a2?a5:a5)):(3'sd1))};
  assign y11 = {{4{(&{{1{(~&p12)}}})}}};
  assign y12 = ({1{{1{$signed((~^b2))}}}}?((p10<=a4)<=(~^a0)):(!(^(a4!=a0))));
  assign y13 = {(|{p5,b4,a5}),(~&{1{a5}})};
  assign y14 = {(5'd19),(+a5)};
  assign y15 = (~^{2{(!((!(~{2{a1}}))^~{1{{1{{4{a4}}}}}}))}});
  assign y16 = ({1{(~{p11,p9})}}>>>{1{(!(3'sd1))}});
  assign y17 = {{(((p16<<<a1)!=(-(a0&p1)))+{(~&{((+b0)&&(p7|a5))})})}};
endmodule
