module expression_00983(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(5'd25));
  localparam [4:0] p1 = ((|((4'd1)?(-4'sd7):(4'sd3)))?((~|(2'd1))?(!(5'sd2)):((4'd2)?(5'sd9):(5'd15))):(((4'sd0)+(2'd2))?((-3'sd0)?(2'd3):(3'd3)):((3'd6)<<(2'd2))));
  localparam [5:0] p2 = ((5'd2 * ((2'd0)^(3'd2)))<<<(((-2'sd0)<<(2'd0))!=((2'd0)==(4'd1))));
  localparam signed [3:0] p3 = {({(-3'sd3)}!={(4'd1)})};
  localparam signed [4:0] p4 = (((5'd24)|(2'sd1))&((5'd22)>=(2'd1)));
  localparam signed [5:0] p5 = (((4'd1)?(2'sd1):(4'sd4))?(^(+((5'd26)?(-5'sd13):(-2'sd0)))):((2'sd0)?(-2'sd1):(3'd6)));
  localparam [3:0] p6 = (3'sd1);
  localparam [4:0] p7 = (((|(~&((-4'sd4)<<(2'd3))))-(-4'sd7))^~(2'sd1));
  localparam [5:0] p8 = (!((((5'd24)?(-5'sd2):(-2'sd1))?((2'd1)?(-4'sd5):(5'd7)):{(2'sd0)})!==({(!(4'd6))}!=(~|((5'd19)<<(5'sd4))))));
  localparam signed [3:0] p9 = (~|((((3'd5)^(4'd1))>>>((2'sd0)==(5'sd5)))<=(((5'sd0)|(4'd0))<(4'd2 * (3'd3)))));
  localparam signed [4:0] p10 = (|((((4'd13)<<<(4'd9))>>(4'sd7))>=(((-3'sd3)|(5'd23))===(~(2'd1)))));
  localparam signed [5:0] p11 = ((-4'sd1)<<<(-2'sd0));
  localparam [3:0] p12 = (4'd2 * ((3'd3)>(3'd7)));
  localparam [4:0] p13 = ((~^(((2'd1)^(5'd14))>>>{2{(3'd3)}}))<<<{1{(-4'sd6)}});
  localparam [5:0] p14 = {{1{{(~{2{(&(-5'sd11))}}),({3{(4'sd5)}}>(~{(5'd12),(-4'sd0),(2'sd0)}))}}}};
  localparam signed [3:0] p15 = (5'd21);
  localparam signed [4:0] p16 = (((3'sd0)?(5'd5):(4'sd4))?{4{(4'd2)}}:((3'd1)?(4'sd2):(-4'sd1)));
  localparam signed [5:0] p17 = (5'd19);

  assign y0 = {p15,a3};
  assign y1 = ((~(^(b3==a5)))!==((b0!=b5)!=(b1^b5)));
  assign y2 = {1{((b0^a3)?(-2'sd0):(p0))}};
  assign y3 = (2'd2);
  assign y4 = ({2{(b3?a3:b3)}}?{3{a3}}:{4{p16}});
  assign y5 = (((+(p7||p12))>>>(p1^~p0))&((^(p5^~p14))<(p11!=p15)));
  assign y6 = (-2'sd0);
  assign y7 = ({(p0==p13),(p2<a3),(b0>=p14)}-((4'd0)?{a4,a3}:(p5^b1)));
  assign y8 = {((p4?b4:p13)<<<(p10||p6))};
  assign y9 = (4'd2 * (~(a0^~a0)));
  assign y10 = (4'd14);
  assign y11 = (p2>p12);
  assign y12 = {p1,p3,p5};
  assign y13 = (3'sd1);
  assign y14 = {2{(4'd2 * {a0})}};
  assign y15 = {2{{3{{1{p2}}}}}};
  assign y16 = (((~&(p9?p1:p14))-((b3<=b3)===(a3+b0)))<($unsigned((p16?p8:p10))>>>(p6?p2:p2)));
  assign y17 = {1{((2'd2)?(((-p10)?(!a5):(~|b0))):((4'sd0)&((a5?b2:p10))))}};
endmodule
