module expression_00853(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+(~|((4'sd1)>>>(4'd15))))|(~(~|{(4'd15)})));
  localparam [4:0] p1 = {(~|(-2'sd0)),((-5'sd0)?(4'd6):(5'd4)),{(4'd4),(5'd10),(3'sd3)}};
  localparam [5:0] p2 = {({(2'd2),(4'sd7),(2'sd1)}?((-4'sd4)?(4'd11):(-4'sd6)):{(3'd2),(-3'sd3)}),{((5'sd10)?(-5'sd1):(-4'sd7))}};
  localparam signed [3:0] p3 = ({4{{2{(4'sd4)}}}}!=(|(!(+(6'd2 * (~^((2'd1)^(3'd6))))))));
  localparam signed [4:0] p4 = {(((3'd4)&&(4'd4))+((2'd0)+(-2'sd1))),{4{(3'sd3)}}};
  localparam signed [5:0] p5 = ({((3'd5)?(2'sd1):(4'sd7)),(~|(2'd3)),((2'sd0)||(2'sd1))}==(^{(~((2'd2)&&(3'd5)))}));
  localparam [3:0] p6 = (-(~|(((3'd7)?(2'd0):(2'sd1))?(|(!(!(-4'sd0)))):(~((3'sd3)?(2'sd0):(5'd7))))));
  localparam [4:0] p7 = ((2'd2)?(!(-2'sd1)):{(-4'sd2)});
  localparam [5:0] p8 = (|(2'd2));
  localparam signed [3:0] p9 = {(&((3'd2)?(5'd4):(-2'sd0)))};
  localparam signed [4:0] p10 = (((2'd1)|(5'd12))<<<((2'd2)+(2'd0)));
  localparam signed [5:0] p11 = ((((3'sd1)==(5'd20))^~{4{(-2'sd1)}})^~(((2'd1)>>(4'd7))-(+(3'd4))));
  localparam [3:0] p12 = {4{{{3{(3'd7)}}}}};
  localparam [4:0] p13 = (~&(~&(4'd1)));
  localparam [5:0] p14 = (((-4'sd4)<=(4'sd4))>(-5'sd8));
  localparam signed [3:0] p15 = (|((((2'sd1)>=(-4'sd7))&((3'sd3)&&(2'd2)))<((~(~|(2'sd0)))>((-4'sd3)!=(-3'sd2)))));
  localparam signed [4:0] p16 = (&{2{(5'sd4)}});
  localparam signed [5:0] p17 = (5'd2 * (4'd9));

  assign y0 = (5'd2 * (b0!==a2));
  assign y1 = ((({1{p0}}^~(5'sd2))!=(-3'sd0))-{1{(2'd3)}});
  assign y2 = ((+{{b2,a1,p17},(-5'sd8),(a4?a5:b2)})<{1{((p6?p4:p15)?(|{p17,b0,p3}):{a5,p6,a4})}});
  assign y3 = (4'd5);
  assign y4 = ((a3?p12:p7)?(p6^b5):(p9%a4));
  assign y5 = (2'd0);
  assign y6 = ((-5'sd9)/a5);
  assign y7 = ({(b3!==a4),(p16^~b4)}>>>($unsigned(p3)|{p9}));
  assign y8 = {3{b1}};
  assign y9 = (|(p15>>p1));
  assign y10 = (+(~((~|b1)?{3{a0}}:(~a4))));
  assign y11 = (|p11);
  assign y12 = (((|(a4===b2))<=$signed((b4===b1)))===({{2{a2}}}<<<$signed({3{b4}})));
  assign y13 = (-3'sd3);
  assign y14 = (p3);
  assign y15 = ((-2'sd0)<(+(b2?b0:b1)));
  assign y16 = ((a2|b3)?(~{1{a3}}):{3{p7}});
  assign y17 = $unsigned((!{(|$signed((&(|(+$signed($signed((!(-(-{{p6,p3,p2},{p10,p10},(~&$signed(p17))}))))))))))}));
endmodule
