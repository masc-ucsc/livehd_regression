module expression_00063(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(((4'd3)?(-3'sd3):(4'd5))>>>(|(5'd16)))}};
  localparam [4:0] p1 = {4{(^(3'd7))}};
  localparam [5:0] p2 = (-(~(5'sd8)));
  localparam signed [3:0] p3 = (6'd2 * {3{(2'd0)}});
  localparam signed [4:0] p4 = ((~&{4{(2'sd0)}})&&(((5'd12)&&(4'd10))|{1{((4'd14)!=(4'd6))}}));
  localparam signed [5:0] p5 = ((-(~&(+((-4'sd3)?(-3'sd0):(5'd7)))))?(-3'sd2):((~&(-3'sd2))?((2'd1)!=(3'sd1)):(!(-4'sd0))));
  localparam [3:0] p6 = {1{((+{(2'd2),(4'sd1),(2'd1)})-(~{1{(4'd10)}}))}};
  localparam [4:0] p7 = ((^{3{(2'd3)}})==={2{{4{(-4'sd4)}}}});
  localparam [5:0] p8 = ((4'sd5)?(-3'sd0):(-5'sd3));
  localparam signed [3:0] p9 = ((((4'sd6)>(-2'sd1))&((5'd28)?(2'sd0):(2'd3)))^(((-5'sd5)&(2'd3))/(5'd17)));
  localparam signed [4:0] p10 = {(3'd3),(3'sd3),(4'sd6)};
  localparam signed [5:0] p11 = ({{(-5'sd5),(3'sd0)}}&((2'd2)!=(2'd2)));
  localparam [3:0] p12 = {((2'd1)!=(-4'sd2)),{2{(3'sd1)}},(~|(3'd1))};
  localparam [4:0] p13 = ((((3'sd0)||(4'sd0))>=(~^(2'sd1)))&&(^{4{(5'sd0)}}));
  localparam [5:0] p14 = (({4{(-3'sd2)}}&((4'sd3)>(-4'sd0)))|(3'sd0));
  localparam signed [3:0] p15 = {2{{1{(~^(((3'sd0)<(2'd0))<((2'sd0)<=(5'sd0))))}}}};
  localparam signed [4:0] p16 = {4{(5'sd12)}};
  localparam signed [5:0] p17 = (((3'd5)?(3'sd0):(2'sd0))<=(((3'd5)?(3'd4):(3'sd0))||((3'd3)?(-3'sd0):(5'd11))));

  assign y0 = {4{b1}};
  assign y1 = ($signed({1{($unsigned(((p16<<p12)!=$signed((p3>=p10)))))}})!=$unsigned((~|(~^(-({4{b3}}===(~|{4{a4}})))))));
  assign y2 = {{(p16<<<a4),(a3&a1)},({a1}?(a1?a1:p8):(^a5))};
  assign y3 = ((~p7)<<(p1|p4));
  assign y4 = ({4{b5}}<((p11==p15)||{4{p0}}));
  assign y5 = (((a3>>b3)===(a4?a1:b0))>(a1?b1:b4));
  assign y6 = (-4'sd4);
  assign y7 = ((a5?a2:a5)?(-4'sd6):(b1?a2:b0));
  assign y8 = (((-2'sd0)!==(^b4))<=(3'sd1));
  assign y9 = ((&(b3?a2:b4))?(~(-{2{a0}})):(&{1{(~|a5)}}));
  assign y10 = ((|((a4>=a4)<=(4'd13)))<<(!((+(+b0))!=(-3'sd3))));
  assign y11 = $unsigned(((a1<<a2)^{2{p2}}));
  assign y12 = ({4{{1{a5}}}}-(4'd4));
  assign y13 = (-4'sd4);
  assign y14 = ((~|(p17?p5:p3))?({p12,p5}<<<(p4?p7:p12)):{2{{p0}}});
  assign y15 = {(-3'sd3)};
  assign y16 = (~(+{1{(3'sd2)}}));
  assign y17 = (-3'sd0);
endmodule
