module expression_00228(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd1);
  localparam [4:0] p1 = ({(!(4'd4))}?((5'd30)?(2'd0):(-4'sd6)):{(-3'sd2),(3'sd1)});
  localparam [5:0] p2 = {2{(~^((~(4'd13))&(~|((2'sd0)+(-2'sd1)))))}};
  localparam signed [3:0] p3 = (4'sd1);
  localparam signed [4:0] p4 = {2{{4{{2{(-5'sd9)}}}}}};
  localparam signed [5:0] p5 = {(4'd8)};
  localparam [3:0] p6 = ({3{((4'd15)?(2'd1):(4'd15))}}|(((2'sd1)^(2'd1))?((4'd4)?(-4'sd2):(5'd30)):(~|(-2'sd1))));
  localparam [4:0] p7 = {((-3'sd2)<<<(-2'sd0))};
  localparam [5:0] p8 = {((5'd6)?(2'sd0):(4'd7)),((2'sd1)|(2'd0)),{(-2'sd1),(4'd15)}};
  localparam signed [3:0] p9 = ((4'd0)?(4'd1):(3'sd2));
  localparam signed [4:0] p10 = (4'd13);
  localparam signed [5:0] p11 = (~(^(~|((|(~&(4'd2 * (~^(5'd21)))))!=(((-4'sd5)<(3'sd0))!=(+((2'sd0)>(-4'sd4))))))));
  localparam [3:0] p12 = {2{(5'd2 * {(2'd0),(5'd25),(3'd0)})}};
  localparam [4:0] p13 = (|({((-5'sd6)&(3'sd2)),(~^(3'sd1)),((5'sd11)?(4'sd6):(2'sd0))}^(((2'd0)<=(5'd18))?(5'd2 * (2'd2)):(|(2'sd1)))));
  localparam [5:0] p14 = ((4'd14)&&(5'd1));
  localparam signed [3:0] p15 = ({3{{(2'sd1),(4'd6),(4'sd4)}}}^{{2{(4'sd1)}},(5'd2 * (4'd2)),{(3'sd1),(3'sd1)}});
  localparam signed [4:0] p16 = (5'sd11);
  localparam signed [5:0] p17 = {3{{2{(5'd8)}}}};

  assign y0 = $signed(b4);
  assign y1 = (+((p10?a5:p10)<<<(p7?p1:p8)));
  assign y2 = ((b4<<b3)-(|a2));
  assign y3 = ((a4)===(b0==a2));
  assign y4 = ((a0>=p10)!={4{a2}});
  assign y5 = {((p12^~p3)+(p2>>p9)),((p7>>>b0)&&(a1>=a0))};
  assign y6 = (&(~(p11>=p6)));
  assign y7 = ($signed($unsigned(a4)));
  assign y8 = ((4'd15)<{(4'sd6)});
  assign y9 = ((^(p11^~p6))<<((+b0)<<<(p8)));
  assign y10 = ((p1?p10:b1)?(b1?b3:a5):(b0<<<a3));
  assign y11 = ((b5|a2)%a4);
  assign y12 = (((a3?b2:b4)?(~b4):(3'd7))?((-a3)?(5'd5):(-a5)):(5'd30));
  assign y13 = (((~|(b0>=a3))&&(&(!(~|a4))))>(~|(~&((~&(|p16))&(~^(!p3))))));
  assign y14 = ((5'd3)<(~(!(~|{4{(p2?b4:p9)}}))));
  assign y15 = {(~&(~|(b5===b4))),(^{(p4&&a0)}),((p16||b4)!=(|p9))};
  assign y16 = {(p0?p3:p10),(p1^~p14)};
  assign y17 = ((-4'sd2)!==((b1===b2)?(b1+a4):(b2?b1:a1)));
endmodule
