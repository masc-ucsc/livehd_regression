module expression_00443(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((((4'sd1)^~(3'd0))<=(6'd2 * (3'd3)))>>>({(4'd2),(3'd6),(4'd12)}?((-4'sd1)?(4'd11):(2'd0)):{(5'd12),(2'd1),(5'sd12)}))};
  localparam [4:0] p1 = ((4'd2)?(-3'sd1):(4'sd5));
  localparam [5:0] p2 = (-3'sd1);
  localparam signed [3:0] p3 = (6'd2 * (4'd4));
  localparam signed [4:0] p4 = (((-3'sd2)|(-2'sd1))<<((2'd1)>>>(4'd10)));
  localparam signed [5:0] p5 = (((-2'sd1)!=(4'd15))?((5'd12)?(-5'sd13):(-4'sd2)):((2'sd1)^(4'sd2)));
  localparam [3:0] p6 = (((5'sd14)?(2'd1):(-2'sd1))<=((3'sd3)/(2'sd1)));
  localparam [4:0] p7 = (&((((3'd4)^~(4'd7))==((5'sd0)?(5'd19):(3'd0)))==((5'd12)?(2'd3):(-5'sd1))));
  localparam [5:0] p8 = ((((-4'sd3)==(-5'sd4))||{(-4'sd4),(5'sd7),(-3'sd0)})==(((5'd8)?(2'd3):(-5'sd15))+((3'd6)^~(3'd6))));
  localparam signed [3:0] p9 = ((5'd22)?(5'sd4):(4'd11));
  localparam signed [4:0] p10 = (~^{(2'sd1),(-5'sd15)});
  localparam signed [5:0] p11 = ((3'd1)?(3'd5):(5'd26));
  localparam [3:0] p12 = (&(&{4{(2'd2)}}));
  localparam [4:0] p13 = (~&(((|(-2'sd0))?(|(3'd1)):((-4'sd3)<=(-3'sd2)))<<<({(4'd2),(2'd1)}?(4'd15):(-5'sd7))));
  localparam [5:0] p14 = (4'd8);
  localparam signed [3:0] p15 = ((5'd18)>>((5'd29)?(2'sd1):(-3'sd0)));
  localparam signed [4:0] p16 = {{{3{(-4'sd0)}}}};
  localparam signed [5:0] p17 = {(({(4'd13)}==((5'd27)&&(5'd13)))<=(3'sd3)),(((4'd10)?(-3'sd0):(3'd6))?((2'sd1)?(4'd15):(-4'sd4)):((5'd2)?(3'd4):(5'sd2)))};

  assign y0 = {$signed((({{a4,b0,a2},{p4,a4},(p12+b2)})=={($unsigned((5'd1))),{p13,a0,b5}}))};
  assign y1 = (|((a2>=p9)+(p3<<<p15)));
  assign y2 = $signed(((a5?a4:a3)===(a1?a0:b2)));
  assign y3 = $unsigned($signed(($unsigned($signed(p10)))));
  assign y4 = {$signed((p11&&p7))};
  assign y5 = $signed((a3^a1));
  assign y6 = ((&((~|p15)?(a0&&p2):(p17?p5:b3)))>>>{1{{2{(|(p3?p5:p2))}}}});
  assign y7 = (({{p16,p10,p7},(p11>=p16)})||(((p10&&p1)&&(p8-p6))==((b4!==b0)>=(p0<=p6))));
  assign y8 = ({$unsigned({2{((p9+p6)^(p17^~p6))}})}<={2{((p2==p17)==(p13&p12))}});
  assign y9 = (p5?p0:p0);
  assign y10 = (~|(~p13));
  assign y11 = {$unsigned((+(^(~^(-{(|a3),{p7}}))))),(&$signed(({{b4,b2,p1},(~b2),(~a2)})))};
  assign y12 = (!(a0?a4:p10));
  assign y13 = ($signed($unsigned(b2))?$signed($unsigned(p4)):(5'd2 * b1));
  assign y14 = {2{(5'd2 * (a0-a1))}};
  assign y15 = ((a1&&b3)^~(3'd2));
  assign y16 = {4{(-5'sd2)}};
  assign y17 = (|{3{{1{(b0||p5)}}}});
endmodule
