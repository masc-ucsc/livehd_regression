module expression_00755(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-3'sd2)?(2'sd0):(4'd6))?((3'd0)?(4'sd5):(4'sd6)):((5'd2)?(2'd1):(3'sd3)));
  localparam [4:0] p1 = {4{({2{(5'sd5)}}<<{2{(3'd6)}})}};
  localparam [5:0] p2 = {2{(4'd5)}};
  localparam signed [3:0] p3 = (({(4'sd4),(2'sd1),(4'd8)}||((-4'sd1)?(3'sd1):(-2'sd0)))?((2'd3)?(3'd1):(3'd5)):(6'd2 * {(5'd12)}));
  localparam signed [4:0] p4 = ({4{(4'sd0)}}<={2{((2'sd0)-(2'sd0))}});
  localparam signed [5:0] p5 = ((~|(-4'sd0))>>{3{(4'd9)}});
  localparam [3:0] p6 = ((6'd2 * {1{{3{(2'd3)}}}})>>(((3'd1)|(3'd1))<<<((-2'sd1)?(3'd5):(3'sd1))));
  localparam [4:0] p7 = ((((5'd15)<<<(3'd2))^((3'sd1)>(4'sd3)))<<<(((3'd4)===(-3'sd0))>>>((4'd1)||(5'd9))));
  localparam [5:0] p8 = ((4'd5)?(-4'sd1):((2'd3)?(2'd3):(5'sd6)));
  localparam signed [3:0] p9 = ((2'sd0)?(4'd1):(-3'sd3));
  localparam signed [4:0] p10 = {(((2'd1)?(2'd3):(-5'sd4))?((4'd5)?(-2'sd0):(2'sd0)):((2'sd1)?(2'd0):(3'd7)))};
  localparam signed [5:0] p11 = {4{(5'sd14)}};
  localparam [3:0] p12 = ((|(~((3'd3)?(5'sd14):(3'd4))))<<<((&(-4'sd4))?((2'sd1)%(-4'sd5)):((2'd2)<(4'sd6))));
  localparam [4:0] p13 = (^(3'd1));
  localparam [5:0] p14 = (({((-5'sd10)>(4'd10))}!==(!{(3'sd3),(2'd1)}))|(~^(&(((4'd6)!==(-5'sd1))||((3'sd3)&&(2'd2))))));
  localparam signed [3:0] p15 = (((~|((2'sd1)!==(5'd11)))+(|((5'sd2)==(2'd2))))>>>((~|(!(-3'sd3)))===((4'd11)>>(3'd6))));
  localparam signed [4:0] p16 = ((((4'd5)!=(2'd3))?((5'd21)?(-5'sd14):(2'd1)):((4'd6)?(2'sd1):(3'sd0)))?(5'sd14):(((-5'sd4)/(2'd3))?(5'd11):((5'sd3)?(2'd1):(5'd3))));
  localparam signed [5:0] p17 = (&(~(-(&(2'd2)))));

  assign y0 = {((b5<<<p13)&&(b3<<p14))};
  assign y1 = (((p2?a2:b1)?(~p10):(~^a3))?((|(3'sd0))/p8):(~&(&(a3?p5:p15))));
  assign y2 = {4{{4{p9}}}};
  assign y3 = (4'd5);
  assign y4 = {4{p17}};
  assign y5 = (~&((~((!p1)==(b2!=b1)))>>>(|$signed({(~&b5),(a5)}))));
  assign y6 = (((p9%p17)-$signed(p6))>>(-5'sd10));
  assign y7 = ((((p13?p5:p12)>>>(p9?p14:p0))?((&$unsigned(p3))<((p12/p11))):((a3^~p4)<=(a1>>>a5))));
  assign y8 = (2'sd1);
  assign y9 = ({4{{4{a0}}}}?({4{b4}}^~(a5===b5)):$signed(((~|p15)!=(~|b1))));
  assign y10 = $signed((((~&p7)||(p10^p13))&&{4{p6}}));
  assign y11 = {{2{p6}},{a3,a4,a4},{2{p3}}};
  assign y12 = (!((b1?b1:b1)!==(b2?a0:a5)));
  assign y13 = (2'sd0);
  assign y14 = (+({1{(5'sd3)}}?(-(3'd1)):(a3?a1:b0)));
  assign y15 = {({1{a1}}<<(p1))};
  assign y16 = {4{(b4-a5)}};
  assign y17 = (~|(|(!((~&(a5<<p9))>>(~^(a0<=a5))))));
endmodule
