module expression_00949(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(!(-{(-(-3'sd3)),(^(3'd3)),((5'd7)?(3'sd0):(3'd1))})),(^(-({(3'sd0)}?(+(2'd3)):{(5'd17),(2'sd1),(5'sd6)})))};
  localparam [4:0] p1 = ((((5'd6)||(5'sd15))-((-3'sd1)?(2'sd0):(4'd9)))-(((4'd14)&&(4'd7))&((3'd4)?(5'd28):(-3'sd3))));
  localparam [5:0] p2 = (-3'sd3);
  localparam signed [3:0] p3 = (((!(-2'sd0))<(&(4'sd3)))?(~|((5'sd6)<=(5'd28))):(((4'sd3)/(-2'sd1))-(!(4'd4))));
  localparam signed [4:0] p4 = {4{(3'd6)}};
  localparam signed [5:0] p5 = ((6'd2 * ((4'd7)?(2'd0):(3'd1)))?((~|(5'd25))^(5'd2 * (2'd3))):((|(-3'sd2))!=(^(2'd0))));
  localparam [3:0] p6 = ((((2'd2)?(2'sd0):(-2'sd1))===((4'd3)==(5'd2)))&&(((5'd4)?(2'd3):(-5'sd7))?((-5'sd7)/(-2'sd0)):((5'd24)+(2'd0))));
  localparam [4:0] p7 = (-{4{(((-4'sd5)!=(3'sd3))===(|(2'sd1)))}});
  localparam [5:0] p8 = ((((4'd3)?(3'd0):(-3'sd0))===((4'd4)-(-3'sd0)))||((4'sd6)?(3'sd2):(2'd1)));
  localparam signed [3:0] p9 = (~&((((4'd3)<=(2'd3))<<<(~|(-3'sd3)))&(!((2'd2)?(5'd9):(5'd20)))));
  localparam signed [4:0] p10 = ((2'sd1)&(3'sd0));
  localparam signed [5:0] p11 = {4{(^(-(+(3'sd1))))}};
  localparam [3:0] p12 = {{{(2'd3)},((-3'sd0)!=(2'd2))},(((5'd20)==(2'sd0))>((-3'sd2)^(3'd0))),(((2'd3)!==(4'd3))^((4'd14)+(2'sd0)))};
  localparam [4:0] p13 = (5'd8);
  localparam [5:0] p14 = {(&(^(|(^((5'd3)+(2'd1))))))};
  localparam signed [3:0] p15 = ((-4'sd3)?(-2'sd0):((2'sd0)?(5'd26):(-2'sd0)));
  localparam signed [4:0] p16 = (5'd4);
  localparam signed [5:0] p17 = ((^(((5'd9)?(-5'sd13):(5'd10))!==(&(-5'sd0))))===(!((&(-4'sd3))-{1{(2'd2)}})));

  assign y0 = ($unsigned(((a0!==a4)||$unsigned($signed(a0))))||(((5'd2 * a0)!==(a4^b1))));
  assign y1 = ((p7<p17)|(3'sd3));
  assign y2 = (-5'sd4);
  assign y3 = (|(|(&(-3'sd0))));
  assign y4 = $signed((!({(+((2'd1))),$unsigned((&(^a4)))}&((~|(~|$signed(b5)))&&(~&(a4<<<p6))))));
  assign y5 = (-3'sd1);
  assign y6 = (~|{4{{1{(~^(a3===b5))}}}});
  assign y7 = ({4{(-4'sd3)}}>={3{(a0>=p16)}});
  assign y8 = (2'd3);
  assign y9 = ((-(a5?b4:p16))?{1{(a3===a3)}}:{(a0!=b5)});
  assign y10 = (4'd10);
  assign y11 = {$signed({{{a5}}}),{$signed(p17),$unsigned(b1)},{$signed(p14),{a0}}};
  assign y12 = (((p6!=p2)>>>(p3<=b3))<<<((p15<p17)<(b3<b5)));
  assign y13 = ({2{(|(p3==p7))}}|(6'd2 * (^{2{p12}})));
  assign y14 = (~({(~|{{b5,a5},(a2!=b5),(p8&&a1)})}<<<{(~&(~|p3)),(~^{a5})}));
  assign y15 = ((({2{p1}}&&(b0?p13:p8))^((~&p14)<=(~|a1)))==(!{3{(!p5)}}));
  assign y16 = (~(!{(^(((~|p2)&(~&a2))|(+{a2,a5,b1})))}));
  assign y17 = (^(!(2'sd1)));
endmodule
