module expression_00068(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{1{{2{(2'd3)}}}}};
  localparam [4:0] p1 = ((-(^((5'd3)||(-2'sd1))))===((~(5'sd13))>(!(2'd1))));
  localparam [5:0] p2 = {{(3'd4),(2'sd1)},(~&(5'sd11)),(~(5'd29))};
  localparam signed [3:0] p3 = (6'd2 * ((2'd0)?(2'd1):(4'd5)));
  localparam signed [4:0] p4 = ((((3'sd1)?(-4'sd4):(-2'sd0))?((-5'sd14)==(-3'sd2)):{3{(2'd3)}})>={(+(-3'sd0)),((-3'sd0)>(3'd1)),(~&(-3'sd2))});
  localparam signed [5:0] p5 = ((^{(~(2'd1)),(~(-5'sd5))})||(|{3{(3'sd3)}}));
  localparam [3:0] p6 = (((3'd4)>={(4'd10),(-5'sd15),(-5'sd14)})^~{{2{((2'sd0)<<<(5'sd0))}}});
  localparam [4:0] p7 = (~{1{(-{4{{1{((5'd14)?(3'sd3):(2'd0))}}}})}});
  localparam [5:0] p8 = (~|((~|(~|(5'd14)))!=((2'd1)>=(4'd3))));
  localparam signed [3:0] p9 = (-(~&{1{{3{(~(4'd10))}}}}));
  localparam signed [4:0] p10 = (-((((4'd6)>=(4'sd7))|(|{4{(-4'sd7)}}))>>>(((5'd0)&(4'd5))==((-4'sd7)<(3'd2)))));
  localparam signed [5:0] p11 = (((3'sd1)^~(-2'sd1))/(-2'sd1));
  localparam [3:0] p12 = {(((5'd28)?(-2'sd0):(3'd1))-((5'sd2)?(-5'sd12):(5'sd3))),((5'd2 * (2'd2))>>>(~&(4'sd1))),(~&((5'd21)?(-2'sd0):(2'd3)))};
  localparam [4:0] p13 = ((2'sd1)^~(-2'sd0));
  localparam [5:0] p14 = (-(~((!((+(-2'sd1))>=((4'd6)<<(2'sd1))))==(~|((|(-3'sd3))&((5'sd6)&(2'd3)))))));
  localparam signed [3:0] p15 = {3{(~|(|{4{(3'd0)}}))}};
  localparam signed [4:0] p16 = ((|((5'sd9)==(-4'sd1)))%(3'd5));
  localparam signed [5:0] p17 = ((((5'd29)<=(4'sd6))-{2{(4'd7)}})-(~^((-5'sd3)>>>(4'sd1))));

  assign y0 = (((a2===a1)<<{(b5)})<=((!((&b4)|(~&b3)))));
  assign y1 = $signed(($signed((((p8)?(-a4):(|b5))?(-2'sd1):(&(~(+(~&b3))))))));
  assign y2 = (&(-{b3}));
  assign y3 = {(+(~{4{p0}})),(4'd8)};
  assign y4 = $unsigned($signed(((~|(^($signed((-a3))|(~^(b0?b2:b0)))))^$signed(((b1?b4:p5)?(~a0):(a0?a2:a0))))));
  assign y5 = ((a0>>>b1)!==$signed((a0)));
  assign y6 = {((p17+p7)?{p11}:(a5?b5:p13)),$unsigned(((b3^b3)===(b3?b5:a5)))};
  assign y7 = $unsigned(((6'd2 * p14)));
  assign y8 = ((!{3{{3{a1}}}})?(^((b1>>b3)?(b0?a0:b3):(a4?p4:a2))):($unsigned({4{b5}})));
  assign y9 = ((-(p14>p13))|{4{p1}});
  assign y10 = (|(({3{p16}}?(p6?p15:a5):(p3?p2:p12))?{2{(p13&p4)}}:((p15>>p15)>>>(p16^~b4))));
  assign y11 = ({b0,p0,p8}||{p1,p8,a2});
  assign y12 = ((b3>>>a3)&$signed(a0));
  assign y13 = ((|(&{2{a1}}))^(&(b4?a2:b1)));
  assign y14 = (4'sd0);
  assign y15 = ({4{b0}}=={2{b3}});
  assign y16 = ((p9|a5)&(5'd2 * p2));
  assign y17 = {4{({4{a1}}-(&b5))}};
endmodule
