module expression_00255(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-3'sd0)?(2'd1):(-5'sd10))+((5'd2 * (4'd0))>=((4'd8)>(2'sd1))));
  localparam [4:0] p1 = {(4'd1),(4'd11),(3'sd0)};
  localparam [5:0] p2 = {1{{2{{3{(5'd14)}}}}}};
  localparam signed [3:0] p3 = {{((5'sd1)?(2'd3):(4'sd4))},((2'sd0)&&(4'sd4))};
  localparam signed [4:0] p4 = ({2{(4'sd0)}}?({4{(-4'sd7)}}>=((2'd2)&(-2'sd1))):(5'd10));
  localparam signed [5:0] p5 = ((-4'sd7)<(5'd18));
  localparam [3:0] p6 = ((|(5'd10))?(+(+(~&(5'sd9)))):((4'd13)?(5'sd1):(2'd0)));
  localparam [4:0] p7 = (4'd15);
  localparam [5:0] p8 = (({2{(-5'sd12)}}^{4{(4'sd5)}})===(((-3'sd2)===(4'd4))&{4{(-3'sd1)}}));
  localparam signed [3:0] p9 = (((3'd0)>(-5'sd13))?(-5'sd12):((-3'sd0)||(-4'sd1)));
  localparam signed [4:0] p10 = (-(~^((5'sd6)||(5'd21))));
  localparam signed [5:0] p11 = (~^({(-2'sd0)}?{(3'sd1),(4'sd6),(4'd4)}:((3'sd0)?(4'd3):(5'd6))));
  localparam [3:0] p12 = ({4{((2'd2)>(-2'sd1))}}!=(~{{2{(2'd0)}},{(2'sd0),(5'd21),(3'sd2)}}));
  localparam [4:0] p13 = {(^((-4'sd6)<<<(4'd3))),{{(3'd4),(-5'sd8)}}};
  localparam [5:0] p14 = ((4'd14)?(4'd0):((4'd13)?((-3'sd1)|(4'd9)):((2'd2)&(-5'sd7))));
  localparam signed [3:0] p15 = ((((5'd7)==(5'd26))?{(5'd15)}:((2'd2)|(5'd21)))||(((2'd0)<(3'sd1))=={(3'd7)}));
  localparam signed [4:0] p16 = (5'sd1);
  localparam signed [5:0] p17 = (5'd9);

  assign y0 = (5'd30);
  assign y1 = (4'd10);
  assign y2 = (5'd2 * (a0?b0:p12));
  assign y3 = (5'd15);
  assign y4 = (((-5'sd12)^((5'd2 * a0)<<<(-5'sd4)))>((a0>=b0)?(p17?p7:a3):(b5!=a2)));
  assign y5 = $unsigned(({{p13,p16,p9},{3{p0}}}>>>((p3?p1:p4)?{p13,p13}:(p14<<<p1))));
  assign y6 = ({(b2^~a1)}?(^{p10,p0,p2}):{p15,p1,p2});
  assign y7 = ((($signed(a1)<{4{a2}})));
  assign y8 = ({(a2>>>a4)}?{a5,b1}:(2'd1));
  assign y9 = (5'd20);
  assign y10 = {3{(a0+a0)}};
  assign y11 = $unsigned($signed({4{{3{b3}}}}));
  assign y12 = ($signed((a3===a1))-(6'd2 * p6));
  assign y13 = ({{(b4&b3)},({b5,a2})}||$signed({(({$signed($signed(a5))}))}));
  assign y14 = {{1{(~^{3{p13}})}},((-a2)&&{2{a3}}),{4{p11}}};
  assign y15 = ({{{p6,p0}},(6'd2 * (5'd9))}||{({4{p13}}<={a3,p1}),((4'd3)^{3{p12}})});
  assign y16 = (({2{(p6-b0)}}&((b3<<b5)>=$signed(p17)))|{1{((p3>=p17)+((b2===b4)))}});
  assign y17 = ((b3?a5:a4)!=((a2<<p9)^~(p15<<<a1)));
endmodule
