module expression_00139(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{(((-4'sd3)?(2'd2):(5'd17))?{3{(4'd13)}}:((3'd0)?(3'sd2):(3'd2))),(~^{2{((-4'sd0)|(5'd7))}})});
  localparam [4:0] p1 = (((!(5'sd6))?((4'sd0)>(5'd14)):(~(2'd0)))?(~|((~(-3'sd0))+(+(-5'sd10)))):((|(2'd2))!==((5'd15)?(3'd1):(4'sd0))));
  localparam [5:0] p2 = {4{((2'd0)===(3'd2))}};
  localparam signed [3:0] p3 = (({(-3'sd2),(5'sd5),(2'd3)}||(|(4'd7)))<<<(((-3'sd2)|(3'd4))==={(-5'sd4),(-2'sd1),(5'sd14)}));
  localparam signed [4:0] p4 = {({(2'sd0),(-2'sd0),(4'd12)}<{(4'd1),(2'd1),(4'd10)})};
  localparam signed [5:0] p5 = {((2'd2)===(2'd3)),((3'd0)<=(-3'sd2))};
  localparam [3:0] p6 = (5'd15);
  localparam [4:0] p7 = ((-(&(-4'sd4)))<=((5'd24)<=(4'd3)));
  localparam [5:0] p8 = ((~|(~^(-3'sd3)))?(2'sd0):(|((-2'sd1)>(5'd19))));
  localparam signed [3:0] p9 = {{((~((-4'sd4)<(5'sd15)))===(|(+(5'd11))))},((|((-3'sd2)|(-5'sd2)))-(6'd2 * (6'd2 * (2'd2))))};
  localparam signed [4:0] p10 = (6'd2 * (3'd0));
  localparam signed [5:0] p11 = {2{(2'd2)}};
  localparam [3:0] p12 = ({(2'd3),(-2'sd0),(-2'sd1)}?(5'd2 * (5'd20)):(3'd7));
  localparam [4:0] p13 = (^({3{(5'd17)}}?{((-3'sd2)+(-5'sd9)),((4'd2)===(-3'sd1))}:{4{(-2'sd1)}}));
  localparam [5:0] p14 = ((~{((2'd0)<<(5'd12)),(~^(-3'sd1)),{(3'd5),(-5'sd14),(5'sd12)}})&({1{((4'd14)>>>(4'sd6))}}<{3{(5'd9)}}));
  localparam signed [3:0] p15 = {(4'd12)};
  localparam signed [4:0] p16 = {{(+{(-3'sd0),(-4'sd6),(-2'sd1)})},({(3'd3),(-5'sd15)}+((4'd10)>>(4'd6)))};
  localparam signed [5:0] p17 = ({4{(5'd26)}}?{{(3'd0),(4'd2)},((-5'sd1)>>(-3'sd2)),((3'd4)<<(-2'sd0))}:{2{((2'd1)>(4'd6))}});

  assign y0 = ((!((~&(p4&&a0))^~(!$unsigned(b2))))<=(!((^((+a1)&&$signed(a4))))));
  assign y1 = (2'sd1);
  assign y2 = ({1{(~(4'd2 * p13))}}|(^{4{p13}}));
  assign y3 = (4'd9);
  assign y4 = $signed((-(2'd1)));
  assign y5 = ((4'sd1)?((p9?p5:p6)?(-5'sd9):(b2?a2:a0)):((p16?a3:a1)/p5));
  assign y6 = {1{(2'sd0)}};
  assign y7 = (~|(5'sd6));
  assign y8 = (+$signed($unsigned(a2)));
  assign y9 = ({p17,p0,b1}&{1{(-3'sd0)}});
  assign y10 = $unsigned((4'sd6));
  assign y11 = {3{{2{(&{4{a5}})}}}};
  assign y12 = {2{{2{(-2'sd1)}}}};
  assign y13 = $signed($unsigned(((a0?p14:p17)^(a2?p3:p0))));
  assign y14 = $unsigned((a3>>>b3));
  assign y15 = ({3{p17}}+{1{{2{b4}}}});
  assign y16 = {(+{(-4'sd2),((+p14)<<<(~^b4)),(+((a2===a3)^(~&p15)))})};
  assign y17 = (((|p0)<<<(b5?p16:p8))?(+((~|b1)>>{b0,a3})):({4{p12}}?(&p17):(b2?a4:b4)));
endmodule
