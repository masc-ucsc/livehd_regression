module expression_00590(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!{3{((3'sd2)?(4'd8):(5'd5))}});
  localparam [4:0] p1 = (^{4{(6'd2 * ((4'd0)&(2'd3)))}});
  localparam [5:0] p2 = (4'd2 * ((4'd12)?(5'd14):(2'd0)));
  localparam signed [3:0] p3 = ((((-4'sd7)!==(3'sd2))-((4'sd3)===(-2'sd0)))?((5'd2 * (4'd12))&((4'sd1)<(4'sd0))):(((3'd6)?(-5'sd7):(5'd9))<<((-2'sd1)^~(3'd1))));
  localparam signed [4:0] p4 = {{(-4'sd6),((3'd7)&&(3'sd0)),{2{(2'sd1)}}},(6'd2 * (~^{(4'd10),(5'd26)}))};
  localparam signed [5:0] p5 = (^(|(&(((-4'sd3)<<<(4'sd5))?{1{(!(4'd8))}}:{4{(-5'sd1)}}))));
  localparam [3:0] p6 = (^{((-3'sd0)?(5'd0):(2'sd0)),(~(5'd21))});
  localparam [4:0] p7 = ((~^{2{{4{(-4'sd6)}}}})||((5'd2 * (5'd27))>>(|((4'd11)!==(-2'sd0)))));
  localparam [5:0] p8 = {2{{(5'd2),(-5'sd0)}}};
  localparam signed [3:0] p9 = ((((2'd1)<<(3'd7))<<<((4'sd7)>>(4'd13)))?({(-5'sd3),(5'sd13)}!=((3'd7)||(-4'sd0))):(((2'sd1)^(-2'sd0))?((2'd3)<(3'sd1)):((5'd10)?(-4'sd4):(3'd5))));
  localparam signed [4:0] p10 = ({(4'd7),(-2'sd0)}===((-5'sd15)<=(2'd0)));
  localparam signed [5:0] p11 = ((2'sd0)+(2'd3));
  localparam [3:0] p12 = (~((-(|(-2'sd0)))?((-5'sd14)?(5'sd6):(2'sd1)):(|(~(3'd0)))));
  localparam [4:0] p13 = ((((3'd6)?(-2'sd0):(2'sd0))?{3{(-5'sd11)}}:((3'd3)^~(3'd2)))+(((-5'sd15)>=(3'd3))-((3'sd1)!=(5'sd13))));
  localparam [5:0] p14 = (6'd2 * ((5'd5)?(2'd0):(3'd0)));
  localparam signed [3:0] p15 = (2'd0);
  localparam signed [4:0] p16 = ((2'sd1)===(-3'sd2));
  localparam signed [5:0] p17 = (~^{(((3'sd0)==(2'd0))&&((2'd3)&&(3'd5))),{(!(((3'd7)-(5'd26))-(~^(3'sd2))))}});

  assign y0 = ((+(a4===b4))?{3{a5}}:(&(a2>a5)));
  assign y1 = {(~|($unsigned((5'd22)))),(~|{$unsigned((&b4)),(3'sd2)}),(~(4'sd1))};
  assign y2 = (|$unsigned((~|(5'sd10))));
  assign y3 = $signed($unsigned({({{a1,b4,b3},(a4>>>b0)}===(((a5|a5)))),{$unsigned((|p5)),$signed((p4>>p9)),{1{{4{p9}}}}}}));
  assign y4 = (!(((b2>>b4)^(a5!==b0))<<((|b4)&(~b1))));
  assign y5 = {({(b4===a0)}^~(4'd2 * $unsigned(p1))),($signed((b5&p6))^($signed(p3)>=(p11^p15)))};
  assign y6 = ((~&(+(!((p6>>p4)/p14))))?(!((~a5)?(&p12):(~&b1))):(|(|((a5!==b5)===(b0?b1:b1)))));
  assign y7 = (^((~&(p11?p11:p17))?(a4?a2:p1):((p4?p4:p6)&(p5))));
  assign y8 = {4{b5}};
  assign y9 = (&(&((b3?p10:a0)?(p14>>a5):(a1>=b3))));
  assign y10 = ((~(-4'sd6))>>{1{(p8|p3)}});
  assign y11 = (|(-3'sd0));
  assign y12 = {2{({1{((5'd29)&(a0<<<b3))}}<<$signed((6'd2 * $unsigned(b4))))}};
  assign y13 = {{{{b5,a1},(~^p9),(a3>=p17)},(~^((b5-b1)&{p2,b1}))}};
  assign y14 = (((^(~|(p9|a4)))>>(-4'sd4))<((~(b5&b4))!==((!b1)>>>(~^a5))));
  assign y15 = (!(a5?a5:b4));
  assign y16 = {(!(~$signed((|((4'sd4))))))};
  assign y17 = (5'sd14);
endmodule
