module expression_00617(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(3'sd0),(((3'd5)^~(3'sd1))>{(4'd1),(5'd19)})};
  localparam [4:0] p1 = (((-(5'd19))|(~&(5'd27)))?((~|(3'd5))||{(5'd20),(2'd3),(3'sd3)}):(~(((-4'sd7)?(2'd1):(-5'sd6))&&{(2'sd0)})));
  localparam [5:0] p2 = (-2'sd1);
  localparam signed [3:0] p3 = ({1{{3{(5'sd10)}}}}?{2{{3{(5'sd6)}}}}:{4{(5'sd15)}});
  localparam signed [4:0] p4 = (4'd2 * ((4'd14)>(4'd1)));
  localparam signed [5:0] p5 = (((~|(~&(3'd3)))|((-2'sd1)<<(3'd1)))+((5'd4)%(4'sd6)));
  localparam [3:0] p6 = ((~(3'd5))^~{2{(5'sd2)}});
  localparam [4:0] p7 = ((2'd3)<=(4'd0));
  localparam [5:0] p8 = (|{(-4'sd2),(2'sd1),(3'd4)});
  localparam signed [3:0] p9 = (~^(6'd2 * ((2'd2)==(4'd12))));
  localparam signed [4:0] p10 = (~(~|((5'sd1)?(4'd14):(-2'sd0))));
  localparam signed [5:0] p11 = {(~(~^(~|{3{(-(2'd3))}})))};
  localparam [3:0] p12 = ({(((2'sd1)<<(4'sd5))>=((5'd26)<<<(2'sd0)))}&&(((5'd9)==(4'd4))?{(-2'sd1),(4'd15),(3'd3)}:((4'sd3)?(5'sd13):(4'd1))));
  localparam [4:0] p13 = ((2'd0)?(4'd7):(-3'sd3));
  localparam [5:0] p14 = (|(~&(-3'sd1)));
  localparam signed [3:0] p15 = (+{4{((5'sd13)<=(-4'sd6))}});
  localparam signed [4:0] p16 = (~{3{((3'sd1)<<(5'd20))}});
  localparam signed [5:0] p17 = {{((5'd8)?(5'd22):(5'd28)),{(4'd15),(-3'sd2)},((3'd1)?(5'd13):(4'd1))},({(5'd23)}?(~|(3'sd0)):(^(2'sd1))),(((5'd30)?(-4'sd3):(4'd15))?(&(-3'sd3)):(-(-5'sd8)))};

  assign y0 = (4'sd4);
  assign y1 = $signed(((b2?b4:p6)?(!p1):{a5}));
  assign y2 = ((3'd4)<<(((a3^~a2)!==(4'sd3))!==((a4<b5)+(a0-a4))));
  assign y3 = {(p11?p1:a0),{p7,p4}};
  assign y4 = ((a3<a2)>>>(a5>>>a4));
  assign y5 = (3'd5);
  assign y6 = (~(~(^{3{p15}})));
  assign y7 = $unsigned({p8,p3,p2});
  assign y8 = ((&{(!(-$unsigned($unsigned(((p0&b4)||(p16!=p8))))))}));
  assign y9 = (p3^~a4);
  assign y10 = {3{(p5||p13)}};
  assign y11 = ((a1<<<b3)%a1);
  assign y12 = (^{{((|{((b3|a2)>={b0,b5})})|{(~&(+b4)),{b3,a4}})}});
  assign y13 = {({b2,p14,p16}>=(2'sd0)),((4'sd2)|(5'sd3)),{(2'd0)}};
  assign y14 = ($unsigned((~&(~&$signed({3{{1{{2{a1}}}}}})))));
  assign y15 = (+(~^b3));
  assign y16 = ((!{4{(p17||p4)}})>=(~&{(p15^p1),(p7|b3),(4'd3)}));
  assign y17 = (((|(a1||a4))==(!(p3<=b0)))?(~|((p6%p13)&&(a4+b0))):((^b2)?(-b5):(b3<=a2)));
endmodule
