module expression_00479(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(5'd26)}};
  localparam [4:0] p1 = (6'd2 * (!(^(5'd2))));
  localparam [5:0] p2 = (~&(&(!(^(2'd2)))));
  localparam signed [3:0] p3 = (~&((2'd0)+(4'sd0)));
  localparam signed [4:0] p4 = {(3'sd1),(-3'sd3),(4'sd5)};
  localparam signed [5:0] p5 = ((((5'd23)>>(4'd10))?((-5'sd3)!=(2'd3)):((4'sd4)-(-3'sd1)))<(((-2'sd0)?(-5'sd8):(2'sd1))/(-4'sd1)));
  localparam [3:0] p6 = (((4'd10)?(3'd7):(2'sd1))?((4'd9)^(-4'sd7)):((3'd2)<(2'd2)));
  localparam [4:0] p7 = ((!(~^(~|(~&(-4'sd5)))))&(((-2'sd1)<=(3'd2))>(&(~&(4'd3)))));
  localparam [5:0] p8 = (~(~((4'd4)<<<(5'd30))));
  localparam signed [3:0] p9 = ((((-5'sd5)?(-4'sd1):(5'sd12))?((5'd28)?(2'd1):(-3'sd3)):((2'd2)>>>(3'd5)))?({(5'd10)}?(4'sd5):((2'sd0)?(5'sd3):(4'sd2))):((5'sd12)|(4'd15)));
  localparam signed [4:0] p10 = ((-3'sd0)?(3'd7):(-4'sd2));
  localparam signed [5:0] p11 = ({(5'sd1),((5'd1)&(3'd5))}||({(5'd5),(-3'sd2)}<{2{(3'sd2)}}));
  localparam [3:0] p12 = ((4'd10)?(4'd3):(3'd6));
  localparam [4:0] p13 = ((~|((4'sd3)&&(-4'sd3)))*(^(|(-4'sd5))));
  localparam [5:0] p14 = ((4'sd6)?(3'd2):(2'd3));
  localparam signed [3:0] p15 = (&(((3'sd3)&(4'sd4))?((2'd2)<(4'd3)):((-4'sd1)/(-3'sd2))));
  localparam signed [4:0] p16 = {{(((4'd7)?(4'd6):(-4'sd1))?((2'd1)?(3'd4):(4'sd6)):(((-2'sd1)==(-4'sd7))+{(-4'sd3),(3'sd0),(4'sd4)}))}};
  localparam signed [5:0] p17 = ((5'sd1)^~(5'sd10));

  assign y0 = {4{{3{(p11|b2)}}}};
  assign y1 = ((~|(-5'sd10))?(-(3'd1)):(5'd15));
  assign y2 = {(((p12?p6:p10)?$unsigned($unsigned(a3)):(p0>>>p0))&&$unsigned(({p8,p8}?{(5'd2 * p12)}:$unsigned((p7<<p0)))))};
  assign y3 = (4'd9);
  assign y4 = (~(^(({1{p7}}|(~&p7))<<<((a3?p2:a0)?(a5^p0):(p14?b1:p8)))));
  assign y5 = {((p9<<<b2))};
  assign y6 = ((b2?b1:a3)?(2'd1):(a0===a5));
  assign y7 = $unsigned({4{(b2)}});
  assign y8 = (((b0|a2)^(a3^~p0))<<({b4}=={a3}));
  assign y9 = $signed(((b3?b4:a5)?(a0?b1:a1):(a0?b4:a2)));
  assign y10 = {p10,p4,p3};
  assign y11 = ((-((~&(+(&p2)))&&((~|p7)<<<(&p13))))<<<(+(|(~&((+(p1<=p16))-(b5>=b4))))));
  assign y12 = (3'd7);
  assign y13 = ({(~|(a3&&a5)),{a3,a3}}^(((a4?a1:a0))||(a3!==a3)));
  assign y14 = ((2'sd1)?((5'd5)?$signed(a4):(5'd6)):(((p10?p5:p17)?{2{p8}}:(2'd0))));
  assign y15 = {2{{3{(~&(~|p5))}}}};
  assign y16 = (4'd5);
  assign y17 = {((p17^~p6)),{{(a1)}},({a4,p12}==(p8>a0))};
endmodule
