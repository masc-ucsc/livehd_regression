module expression_00667(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd5)^~(-3'sd2))?(5'd30):(6'd2 * (4'd5)));
  localparam [4:0] p1 = (((3'sd2)>>(4'd14))/(-2'sd1));
  localparam [5:0] p2 = ((((5'd9)?(5'd25):(-2'sd0))^~((3'sd3)===(2'sd0)))>={1{((-2'sd1)?((3'd0)^~(2'd3)):(2'd3))}});
  localparam signed [3:0] p3 = (~&((3'd3)+(~&(5'd25))));
  localparam signed [4:0] p4 = (&{1{{(((4'd1)>>>(4'd8))&((2'd1)^(-2'sd0))),(!((~^(5'sd11))<{(-5'sd8),(-3'sd1)})),({3{(2'd0)}}<<((4'sd5)^~(-4'sd0)))}}});
  localparam signed [5:0] p5 = ((-4'sd4)||(2'd2));
  localparam [3:0] p6 = ((^((6'd2 * (5'd0))<=(!(~&(-4'sd3)))))<=(-((^{4{(4'd1)}})^((4'd0)&&(4'd3)))));
  localparam [4:0] p7 = (3'd5);
  localparam [5:0] p8 = (|(|((~|(~|(|(|(3'd6)))))===(((4'd11)>(3'd5))&&((5'd23)!==(5'd15))))));
  localparam signed [3:0] p9 = (~^(3'd1));
  localparam signed [4:0] p10 = {{1{((-5'sd8)+{3{(3'd2)}})}},{(-2'sd0),{(5'd4)}}};
  localparam signed [5:0] p11 = {2{(-3'sd1)}};
  localparam [3:0] p12 = (((5'sd8)&(3'd1))?((4'd12)-(-3'sd1)):((2'd3)?(5'd30):(5'd10)));
  localparam [4:0] p13 = (2'd0);
  localparam [5:0] p14 = {2{((-3'sd2)?(3'd6):(-5'sd10))}};
  localparam signed [3:0] p15 = (((4'sd3)>=(-4'sd0))===((-4'sd0)!=(-5'sd4)));
  localparam signed [4:0] p16 = (-4'sd7);
  localparam signed [5:0] p17 = {1{(2'd0)}};

  assign y0 = {(5'd2 * {p7,b0}),((b5<=p13)&&(a0!==a4))};
  assign y1 = ($unsigned({2{{4{(p0)}}}}));
  assign y2 = (a4-b2);
  assign y3 = (((p3?a4:p8)<<(2'd2))?((p17?p7:p15)?(a0?p1:p9):(3'd3)):((p3^b4)>(p9?p7:p1)));
  assign y4 = ((+(4'sd1))?(4'd5):(a3?b3:p14));
  assign y5 = $unsigned($unsigned($unsigned((^$unsigned((^(~|((b4==p17)>>>{1{p7}}))))))));
  assign y6 = {b1,p13,p16};
  assign y7 = (((p15<<a5))?(b4===a4):(a2?b1:b1));
  assign y8 = (^(((+p5)?(2'd3):{3{a2}})?(-3'sd2):(+{2{{p4,p10}}})));
  assign y9 = ($signed(p15));
  assign y10 = (((+{2{b1}})>{1{(~(-b1))}})==(((b0==a0)||(a2!==a0))>>((a1>a5)>={3{p16}})));
  assign y11 = ((~|(&(~^(!(~{3{a2}})))))?(({2{b4}}>(~(b2?a4:a1)))):{2{(2'd2)}});
  assign y12 = (((a1?b2:p2)?(b1===b4):(a3?p13:p0))==((b4?p17:b2)>=(p6?p7:p10)));
  assign y13 = (p12==p4);
  assign y14 = ((+((a4|p7)*(^(a3<<<a4))))-((~|(a4!=p2))==(p4==b3)));
  assign y15 = (4'd15);
  assign y16 = (~|(((a0!==a3)>{a1})?(a2?a3:a3):(a5?b2:p2)));
  assign y17 = ({2{((b1+b4)===(~&(a4^a5)))}});
endmodule
