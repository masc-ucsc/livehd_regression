module expression_00083(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({3{(2'sd0)}}?{3{(5'sd6)}}:(|{((2'sd0)?(3'd4):(3'sd3))}));
  localparam [4:0] p1 = {(~^({(4'd13),(3'sd0)}?{(5'd18)}:((5'sd0)?(4'sd0):(3'd2)))),(|(!{(4'd8),(2'd1),(4'sd4)}))};
  localparam [5:0] p2 = ({(~^(2'd1))}>>(5'd2 * (2'd0)));
  localparam signed [3:0] p3 = ((5'd4)?(-5'sd4):(3'd7));
  localparam signed [4:0] p4 = ((^((-2'sd0)^(4'sd7)))+{1{(~{4{(3'sd3)}})}});
  localparam signed [5:0] p5 = (+(((!(2'd1))&(~|(2'd2)))!=(((2'd2)>=(3'sd3))===(&(5'sd12)))));
  localparam [3:0] p6 = ({2{(3'd7)}}^~{2{(-3'sd3)}});
  localparam [4:0] p7 = (-5'sd7);
  localparam [5:0] p8 = {2{{4{(5'd26)}}}};
  localparam signed [3:0] p9 = ((+((5'sd7)?(2'sd0):(5'sd9)))>>>(~|((5'sd15)?(3'd6):(-4'sd2))));
  localparam signed [4:0] p10 = (((4'd6)!==(-4'sd6))>>>(-2'sd1));
  localparam signed [5:0] p11 = (&(3'd1));
  localparam [3:0] p12 = ((^(3'd6))!==((~&(4'd15))<=((-4'sd3)?(2'sd1):(3'd2))));
  localparam [4:0] p13 = (((-{1{(5'd28)}})!=={3{(-3'sd1)}})<<<(-3'sd1));
  localparam [5:0] p14 = {2{(5'd2)}};
  localparam signed [3:0] p15 = ((((3'd2)||(-2'sd1))||{(-2'sd1),(4'd13)})&(((3'd5)?(4'd3):(4'd4))||((4'sd5)&(4'd7))));
  localparam signed [4:0] p16 = (~(^(~&({(2'd2),(-2'sd1),(3'sd0)}>>>((2'd0)!==(4'd15))))));
  localparam signed [5:0] p17 = ((~(((3'd4)==(3'd2))>=((-4'sd4)!==(4'sd6))))+{3{((-4'sd5)<=(3'd2))}});

  assign y0 = ((((a5?p16:p8)>(a1>>p1))>=($unsigned(a4)<<(b2>>b3)))-$signed((~&{(5'sd6),(a4===b1),{b5}})));
  assign y1 = (~|(((p11/p7)*$signed((p11)))?($unsigned((^b0))^~(a1<=b5)):((|(+b2))%a2)));
  assign y2 = (^{3{(a5-p8)}});
  assign y3 = ({(p3==a2),(-4'sd2)}?((4'sd4)^~(5'd11)):(!({b4}?(^a5):(~^p9))));
  assign y4 = $signed((((p3?p5:p1)?(~^$signed(p12)):(p13<<<p9))>((~|(p10&&p7))?(p2?p1:p0):(~|(p9&&p3)))));
  assign y5 = (5'd2 * (2'd3));
  assign y6 = (-{4{(-(~(^b4)))}});
  assign y7 = ((-(~&$unsigned(({(a2!==b3),(!(p6>p2))}&((p6>>b5)&&(4'd9)))))));
  assign y8 = ({3{a5}});
  assign y9 = ((((b2^~a5)>>>(a4+b2))>((5'd2 * b1)))&($unsigned({2{p16}})^((b3-b4)+(b3<=b3))));
  assign y10 = ((5'd31)||(((2'd3))>>>(&(~&p4))));
  assign y11 = (p14?p15:p12);
  assign y12 = $unsigned(((b4>=a4)<(p17?p7:b2)));
  assign y13 = ((((a0===b3)!=(p1||p4))&(!(p2^p10)))<(4'd2 * (~^(b1!==a0))));
  assign y14 = {3{{1{$unsigned(p9)}}}};
  assign y15 = (|b0);
  assign y16 = ((5'sd8)?(b0===a3):(b1==p12));
  assign y17 = ((&{(p17<=p4)})?((p14)^~{a2,a5}):{(a4?p4:p3),(|a3)});
endmodule
