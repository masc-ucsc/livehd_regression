module expression_00555(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(((-4'sd3)>(-5'sd11))<<<(5'd27))}};
  localparam [4:0] p1 = {({(-3'sd0),(5'd13),(-4'sd0)}?(-3'sd1):((|(-3'sd1))+((-2'sd1)?(2'd3):(4'd9))))};
  localparam [5:0] p2 = (-3'sd0);
  localparam signed [3:0] p3 = (~&((((-4'sd6)?(4'sd6):(3'sd2))?(^(5'sd7)):(-(5'd9)))>=(|(((4'd15)?(2'd2):(-3'sd1))*((3'd3)>(2'd1))))));
  localparam signed [4:0] p4 = (((-4'sd0)?(3'sd1):(5'd3))<<((-4'sd5)?(2'sd0):(-5'sd12)));
  localparam signed [5:0] p5 = (^({1{(^(5'sd5))}}?((5'd31)!=(5'd10)):((5'd21)!=(3'd2))));
  localparam [3:0] p6 = {(((5'sd3)-(2'd2))<<((-3'sd2)>=(-3'sd2))),{((2'sd1)>(-3'sd0)),(-3'sd2),{(3'sd0),(5'd21),(4'd12)}}};
  localparam [4:0] p7 = ((^((-3'sd1)?(5'd10):(3'd5)))?(4'd13):((5'd30)?(5'd7):(-5'sd11)));
  localparam [5:0] p8 = (~{4{(~^((5'd23)?(2'd0):(2'd2)))}});
  localparam signed [3:0] p9 = {2{{1{((5'sd10)!=(2'd0))}}}};
  localparam signed [4:0] p10 = ((4'd6)||(3'd4));
  localparam signed [5:0] p11 = (^{(3'd7),(-2'sd1)});
  localparam [3:0] p12 = {4{(-2'sd0)}};
  localparam [4:0] p13 = ((5'sd8)?((4'd9)?(3'd1):(2'd1)):{4{(5'd26)}});
  localparam [5:0] p14 = ((-3'sd3)^~(-5'sd5));
  localparam signed [3:0] p15 = ((~|(^(~&(((5'sd8)<<(3'd0))<((5'sd13)>=(4'd3))))))&(((5'd26)&&(-5'sd7))-((-2'sd0)*(5'd15))));
  localparam signed [4:0] p16 = ((3'sd2)?(4'sd1):(5'd2));
  localparam signed [5:0] p17 = (|(-(+(((~|(2'sd1))-{4{(-3'sd0)}})!==(|{4{(-5'sd11)}})))));

  assign y0 = (~(-{4{(6'd2 * p6)}}));
  assign y1 = {4{(2'd1)}};
  assign y2 = (a4<a2);
  assign y3 = (~^$unsigned($signed($unsigned($signed((~&(~&(~|(+((-(~|(b0<<<a3)))))))))))));
  assign y4 = (a0<a3);
  assign y5 = (~{1{{{1{({b5}^~{p8})}}}}});
  assign y6 = ((p11?b0:b4)>(a3?b3:b4));
  assign y7 = ({4{p6}}<<<((a4&&p14)^(4'd2 * p2)));
  assign y8 = (-5'sd12);
  assign y9 = (($signed({(a4<=b5),(p12^~p13)})>>>({(p3==p3)}=={p3,p12,p7})));
  assign y10 = (-(^(2'sd0)));
  assign y11 = (((a5?b1:b4)<=(-(b1?a4:b0)))!=={3{{2{b3}}}});
  assign y12 = ({(2'd2),{p5,p0,p3}}|(2'd1));
  assign y13 = (((b3===a4)===(-a5))>>>{(b5<<a1),(a2>>>a0)});
  assign y14 = ({3{p6}}?(a2?b1:a4):(2'd3));
  assign y15 = (((5'd12)?(+p11):(+a1))?((b0?a3:b2)>>$unsigned({b5,a1,p1})):(+(5'sd5)));
  assign y16 = (!{4{(~^(4'sd2))}});
  assign y17 = {4{(b1>p3)}};
endmodule
