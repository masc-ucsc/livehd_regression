module expression_00351(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(~^(^(2'sd0))),{(&(5'd15))}};
  localparam [4:0] p1 = (~^(!(4'sd4)));
  localparam [5:0] p2 = (((3'sd3)&(2'd0))>>(~&(3'd4)));
  localparam signed [3:0] p3 = {{(5'd11)}};
  localparam signed [4:0] p4 = (({1{(5'd6)}}+((5'd11)||(-5'sd11)))^~{3{(5'sd8)}});
  localparam signed [5:0] p5 = {(2'sd1),(4'd11)};
  localparam [3:0] p6 = {3{{4{(-5'sd0)}}}};
  localparam [4:0] p7 = {1{{1{(^(3'd4))}}}};
  localparam [5:0] p8 = (|{({(3'sd2),(3'd7),(5'd23)}>(~^(5'd5))),{{(-4'sd4),(4'd6),(3'd1)},(&(2'd3))},{(~^(-4'sd4)),((5'd11)===(-4'sd4)),{(5'd18),(2'sd0)}}});
  localparam signed [3:0] p9 = ((((-4'sd0)+(4'd10))==((3'd7)<<<(-2'sd1)))>>>(((2'd1)||(2'sd1))===((4'sd4)>>>(5'd25))));
  localparam signed [4:0] p10 = ((~(3'sd1))!=((-3'sd2)+(~^((4'sd6)>>(5'sd14)))));
  localparam signed [5:0] p11 = ((((2'd2)>(-3'sd0))%(2'd1))>>(((-3'sd0)/(3'sd1))%(3'd0)));
  localparam [3:0] p12 = {3{(((5'd10)&&(5'd21))==={1{(2'd2)}})}};
  localparam [4:0] p13 = (5'd27);
  localparam [5:0] p14 = {((((3'd1)?(4'sd5):(3'd4))?((2'sd1)?(2'd2):(3'd3)):((3'sd2)!=(5'sd3)))||(((4'd0)?(5'd3):(4'd7))?((4'sd7)?(-2'sd0):(4'd15)):((3'd1)&(3'd1))))};
  localparam signed [3:0] p15 = (6'd2 * (~(~(5'd11))));
  localparam signed [4:0] p16 = (((4'd15)!=(-3'sd1))!=(4'd5));
  localparam signed [5:0] p17 = {2{{(4'd1),(2'sd0),(-5'sd10)}}};

  assign y0 = ((((4'd2 * p8)<<<(6'd2 * p13)))<=({p16,p1}>>>(p12^p9)));
  assign y1 = (~|$signed((|(~^(5'sd14)))));
  assign y2 = (~{(p2?p2:a4),{3{p1}},(~a4)});
  assign y3 = ((p16?p7:p17)?{p13,p10,p5}:{p17,p2,p11});
  assign y4 = (~&(((|p10))?(~&(|p10)):(&(~&b4))));
  assign y5 = (3'd7);
  assign y6 = $unsigned({(-{(b3===a2),(!(a4>b4)),(5'd2 * p6)}),({1{($signed((b4==a5))!=(b4||b1))}})});
  assign y7 = ((3'd6)|((&(3'd3))<<((-2'sd1)>>>$signed(p4))));
  assign y8 = $signed(((((4'd2 * $unsigned($signed(b1)))^{((b1<<a3)>>>(p5<<<p0)),((b2>b4)-{b1,a2,a1})}))));
  assign y9 = ((((p6>p2)!=(4'd13))&&(3'd1))!=(5'sd2));
  assign y10 = (3'd7);
  assign y11 = (~($signed(((b3?a0:a5)&(a0===a4)))&&({1{b2}}&&$signed(a0))));
  assign y12 = ((p5||b0)/a1);
  assign y13 = {3{(~&$signed((b3?a0:a2)))}};
  assign y14 = ((2'sd1)>=(((a3<<<b1)===(a5*a1))!==(-3'sd3)));
  assign y15 = (2'sd0);
  assign y16 = $unsigned({{(+($unsigned((p13&&p0))>=(p1|p2))),{((p12<<<a4)>(~{a4,a3,p0}))}}});
  assign y17 = (3'sd3);
endmodule
