module expression_00580(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-((3'sd2)&&(4'd9)))?(-(~(3'sd3))):(~|{2{(4'sd5)}}));
  localparam [4:0] p1 = (((2'sd1)!=(5'd8))<((3'd6)+(5'd27)));
  localparam [5:0] p2 = (+(~&(~(&{2{(-(|{(-3'sd1),(-5'sd13),(-5'sd4)}))}}))));
  localparam signed [3:0] p3 = (&{(&(2'd1)),(2'd2)});
  localparam signed [4:0] p4 = ((5'd2)?((2'sd1)?(5'd14):(4'd11)):((2'sd1)||(-2'sd1)));
  localparam signed [5:0] p5 = (((4'sd4)?(2'd1):(3'd2))?((-2'sd1)<<<(2'd0)):((4'sd4)?(-4'sd3):(3'd7)));
  localparam [3:0] p6 = (-{(5'sd0)});
  localparam [4:0] p7 = (~(+((|(~&(2'd2)))<=((2'd2)&(4'd8)))));
  localparam [5:0] p8 = {(3'd0)};
  localparam signed [3:0] p9 = (~(~^(~((~{(((4'sd6)<<(5'd25))|(~|(4'sd1)))})>>(((4'd11)>(5'd26))!=((-5'sd0)|(-3'sd0)))))));
  localparam signed [4:0] p10 = (~^(5'd16));
  localparam signed [5:0] p11 = (-3'sd2);
  localparam [3:0] p12 = (~^((~&(^(-4'sd2)))?((3'd2)?(4'd1):(5'sd10)):(~&((4'sd6)<<<(-2'sd1)))));
  localparam [4:0] p13 = {((!(4'd9))&&(+(-5'sd12))),(5'sd14)};
  localparam [5:0] p14 = (((4'd5)?(-5'sd0):(3'd7))>>(4'd2 * ((5'd24)?(4'd2):(3'd3))));
  localparam signed [3:0] p15 = (!(((4'd1)?(2'd1):(4'd14))-((4'd15)?(5'd13):(3'sd3))));
  localparam signed [4:0] p16 = (3'd1);
  localparam signed [5:0] p17 = (-{3{((-5'sd10)?(-5'sd14):(-4'sd6))}});

  assign y0 = (~{3{{1{((p16?b3:a4)?(!b4):{2{p10}})}}}});
  assign y1 = (~^($unsigned(((~^b1)&(a4<=b3)))?($unsigned($unsigned(a5))<<(p4>=p7)):((3'd6)|$unsigned((a5?b0:a0)))));
  assign y2 = ({3{(~&(p6^~a5))}}<<<{3{$signed((p5|p15))}});
  assign y3 = (+(a0&b5));
  assign y4 = (-3'sd2);
  assign y5 = (-(3'd5));
  assign y6 = ((&{2{p11}})>=(!(a3<<p14)));
  assign y7 = {(-2'sd0)};
  assign y8 = {1{{2{(&(~&{4{a5}}))}}}};
  assign y9 = {b5,p1};
  assign y10 = ({(a4-p6)}&(5'd31));
  assign y11 = {(+((-{p9,a1})||(~&(a5!=a4)))),((b4|a3)===(b3>>b0)),((6'd2 * b0)<(b1<<<b1))};
  assign y12 = (-$unsigned($unsigned($signed((b4?a0:b1)))));
  assign y13 = {2{{(4'sd1),($signed(a2)?(-5'sd11):{3{b1}})}}};
  assign y14 = (+(((~&(-b4))<<<(p9?p1:p12))<<(|(3'd0))));
  assign y15 = (-(((p14>>>b0)<=(-(a5!=p13)))?(&{1{((!b4)<<<(~p9))}}):{2{(p3==p5)}}));
  assign y16 = (~(({4{b3}}&&{3{p16}})<<((~(&b4))==={2{b5}})));
  assign y17 = ({p16,p3}?(b4|p1):{3{p12}});
endmodule
