module expression_00369(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^{(5'd9)})=={2{(4'd13)}});
  localparam [4:0] p1 = (^((~(((-5'sd9)^(4'd1))?(^(5'sd15)):((4'd2)&(2'd2))))-((~|((4'sd3)?(5'sd7):(5'd31)))>>((3'sd1)<(-5'sd7)))));
  localparam [5:0] p2 = (((-2'sd0)?(3'd7):(2'd0))-(2'sd1));
  localparam signed [3:0] p3 = {3{(-2'sd1)}};
  localparam signed [4:0] p4 = ((4'sd2)!=(3'd3));
  localparam signed [5:0] p5 = ((((2'sd0)?(5'd30):(-4'sd4))===((5'd4)^~(-2'sd0)))-{((5'd11)>(4'sd6)),((-5'sd3)===(2'sd1))});
  localparam [3:0] p6 = {(5'sd14),(4'd7)};
  localparam [4:0] p7 = ({((4'd5)?(3'd4):(-5'sd4))}?{(3'd6),(2'sd1)}:(&((4'd7)?(5'd9):(-2'sd1))));
  localparam [5:0] p8 = (!(-(&(~^(-(((3'sd1)&(5'd22))===(+((-4'sd3)>(-5'sd13)))))))));
  localparam signed [3:0] p9 = (~^(^((^(-3'sd1))<=(~^(!((4'd5)?(-2'sd0):(3'd6)))))));
  localparam signed [4:0] p10 = (((4'd9)<(~&(&(5'd25))))&&(4'sd1));
  localparam signed [5:0] p11 = (({4{(4'd4)}}?{1{((-2'sd0)<<<(5'd5))}}:{1{{2{(2'd0)}}}})&{4{(5'd2 * (4'd12))}});
  localparam [3:0] p12 = {4{(-((-4'sd7)===(2'sd1)))}};
  localparam [4:0] p13 = (6'd2 * ((2'd1)+(5'd8)));
  localparam [5:0] p14 = {{(-2'sd1)},{(4'd9),(5'sd4)},(&(3'sd3))};
  localparam signed [3:0] p15 = (((2'sd0)&(2'sd0))===((3'd5)===(3'd4)));
  localparam signed [4:0] p16 = ((|(-3'sd3))?((4'd10)?(2'd1):(2'd2)):((5'sd3)?(5'sd3):(-4'sd1)));
  localparam signed [5:0] p17 = ((-4'sd1)!==(((5'd28)&(4'sd2))+((5'sd9)-(5'd14))));

  assign y0 = (p2>=p15);
  assign y1 = ((p15?a2:b4)?(2'd2):{b5,p2,p12});
  assign y2 = (4'd8);
  assign y3 = $signed(p10);
  assign y4 = (!(2'd1));
  assign y5 = $signed(((~((+p15)|(p16>p12)))>((p11&p16)==(p15?p16:p1))));
  assign y6 = (4'sd7);
  assign y7 = {(2'd3)};
  assign y8 = ((p7?p10:p4)?(p10?a4:p14):(-2'sd1));
  assign y9 = (~|p7);
  assign y10 = $unsigned({$unsigned($signed({2{a2}})),((b3-a1)<<{b4,b0}),{4{b3}}});
  assign y11 = ((+((5'sd3)?(p16<<<p1):(a3?a5:a1)))|(&({3{a0}}>(|{2{p6}}))));
  assign y12 = (+(!{1{{3{(b2==a2)}}}}));
  assign y13 = (-3'sd2);
  assign y14 = {(+(5'd5)),(~&((|p15)<=(~p17))),$signed({(-4'sd0),{p2}})};
  assign y15 = ((5'd26)<(({b3}>>>$signed(b4))!==(2'd0)));
  assign y16 = (({$signed(p5),(b5!==a0),(p9|b2)})&{3{(b1?p16:a4)}});
  assign y17 = (4'd2 * (p6!=p1));
endmodule
