module expression_00207(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(({4{(-5'sd0)}}&&(+(4'sd7)))<=({(3'sd1)}>{4{(4'd6)}})));
  localparam [4:0] p1 = {{(^(3'd3)),{(2'd3)},(~&(-5'sd12))},(|{(~&(4'd4)),(&(3'd2))}),(~^(^(-{(5'd20)})))};
  localparam [5:0] p2 = ((-5'sd9)^(3'sd1));
  localparam signed [3:0] p3 = (({3{(-5'sd4)}}==(~^((3'sd3)^~(3'd4))))||(-3'sd3));
  localparam signed [4:0] p4 = {(~(2'sd0)),(-(-4'sd6)),{1{(2'd2)}}};
  localparam signed [5:0] p5 = (-{2{{1{(&(3'sd2))}}}});
  localparam [3:0] p6 = (5'd10);
  localparam [4:0] p7 = ((|(5'd7))?((4'd10)?(-5'sd9):(5'sd12)):((4'd2)?(2'd2):(2'd2)));
  localparam [5:0] p8 = (((((-5'sd1)+(2'sd0))>>>(-(3'sd0)))>(((3'd5)%(2'd3))&((5'sd4)|(5'd31))))>>>((((4'd14)>=(5'd24))-((2'd1)/(4'd9)))-(((4'sd5)*(3'd6))^(-(4'd12)))));
  localparam signed [3:0] p9 = (-{1{(^(((5'sd9)>(2'd3))>{(-3'sd2),(2'd2)}))}});
  localparam signed [4:0] p10 = (+{1{(!(~^{4{(4'd13)}}))}});
  localparam signed [5:0] p11 = ((3'sd2)<((5'sd7)===(3'd3)));
  localparam [3:0] p12 = (3'sd3);
  localparam [4:0] p13 = (((5'd1)>>>(5'd6))!=((5'd5)>>(3'd4)));
  localparam [5:0] p14 = (~|(6'd2 * {1{((5'd28)^(2'd3))}}));
  localparam signed [3:0] p15 = (^(~|(~&(3'd6))));
  localparam signed [4:0] p16 = ((-4'sd6)===(5'sd7));
  localparam signed [5:0] p17 = (((-2'sd1)?(4'd14):(2'sd1))?(5'd2 * {1{(4'd11)}}):((2'sd1)?(-4'sd0):(3'd6)));

  assign y0 = (p15?b4:a5);
  assign y1 = ((^(((p1)?(p17):(p12))!=((|b3)?$unsigned(a3):(p7*p7)))));
  assign y2 = ((4'sd6)===(4'd10));
  assign y3 = ({(~&(~&b4)),(a5===a1),(!(-a4))}+{{b1,a4},(~|{b1}),(~(b2<<a5))});
  assign y4 = (~&(~^{((a5<b1)>>(~|(b3-p13))),{(6'd2 * p8),{b0,b0,b5},{a1,a2}},(~&((a4^p14)<=(|b0)))}));
  assign y5 = ((((p14&&a5)-(a0?a5:b3))^~(b4?b3:b2))||(((p12?b0:a5)<(b1<<<a3))!=((b1<<p4)<=(p13?b4:a0))));
  assign y6 = ($signed(((2'sd0)?{b2,a4,a3}:(a2))));
  assign y7 = ((b0>>>a5)+(p0>=p1));
  assign y8 = ((5'sd3)&&(-5'sd0));
  assign y9 = (~|b1);
  assign y10 = (~|(~^((-2'sd0)&(p14%b0))));
  assign y11 = (({1{{p17}}}>={1{(a2>=p5)}})||(~({a5,p4,a1}=={1{{2{a3}}}})));
  assign y12 = $signed(((b5<<<a1)-{a1,a4,p6}));
  assign y13 = ({p5});
  assign y14 = {3{{1{{1{{{2{p4}},{p11,p1},(p11)}}}}}}};
  assign y15 = (~&{2{p5}});
  assign y16 = ((((4'd8)))|$unsigned((3'd0)));
  assign y17 = {{1{$signed(b4)}},{a1,a4},$signed({b2})};
endmodule
