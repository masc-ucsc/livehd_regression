module expression_00311(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd7);
  localparam [4:0] p1 = (((3'sd0)?(-5'sd6):(3'sd0))?(-(^((4'd15)?(4'd15):(5'sd7)))):((4'd2 * (3'd3))<=(3'sd2)));
  localparam [5:0] p2 = (2'd2);
  localparam signed [3:0] p3 = ((^(3'sd0))?(~^(3'd1)):(|(5'sd3)));
  localparam signed [4:0] p4 = (((&(-(5'd22)))<=((-5'sd11)<<(2'd2)))!==(~&(((-4'sd5)&(4'sd7))|(+(4'd2 * (2'd0))))));
  localparam signed [5:0] p5 = ((((2'sd1)?(5'd4):(3'd6))>((4'd0)|(5'sd0)))|(((-2'sd1)?(-3'sd0):(5'd27))-(3'd2)));
  localparam [3:0] p6 = (6'd2 * (2'd1));
  localparam [4:0] p7 = ((5'd1)?(3'd1):(2'sd1));
  localparam [5:0] p8 = ((2'sd0)!==(((5'sd15)!==(3'd4))?((2'sd0)+(5'd3)):((5'd4)?(3'd7):(-5'sd15))));
  localparam signed [3:0] p9 = ((4'd14)>>(((4'sd7)<(5'd19))&((-2'sd1)==(3'd1))));
  localparam signed [4:0] p10 = {((5'd13)?(2'd3):(5'd0)),((5'd3)?(2'sd1):(3'sd3)),((&(3'd2))>={(5'd16),(2'd1),(2'sd0)})};
  localparam signed [5:0] p11 = (((+(5'sd7))?(2'd2):(3'sd1))|{3{{2{(5'sd7)}}}});
  localparam [3:0] p12 = ((-4'sd6)?(4'sd7):(4'd11));
  localparam [4:0] p13 = ((~&((2'd3)?(3'd2):(3'd1)))?(((5'd29)>=(5'd25))&&{(2'd0),(-2'sd1),(2'd2)}):(((-3'sd3)?(2'd0):(2'd0))==((5'd18)<<<(5'sd12))));
  localparam [5:0] p14 = (-2'sd0);
  localparam signed [3:0] p15 = (~|(5'd8));
  localparam signed [4:0] p16 = {((4'd6)?(2'sd0):(4'd4)),((5'd27)?(5'sd8):(2'd3))};
  localparam signed [5:0] p17 = {4{(2'd1)}};

  assign y0 = {1{{a2,b0,a5}}};
  assign y1 = $unsigned(((-4'sd4)&((p5?a0:a4)||$unsigned(a3))));
  assign y2 = (({a3}^(b5|b5))?((b0&&b5)<(b4===b4)):(~(^(a0^~a5))));
  assign y3 = $unsigned({{{3{p13}},(p2!=p9),(p10)},{$signed(p11),(p15^~p10),$signed(p8)}});
  assign y4 = (-2'sd0);
  assign y5 = ({3{p5}}?(!(p14^p7)):(~(p12<=b4)));
  assign y6 = (({b4}<=(a5))^~((b1<<a2)?(a3<b5):(~^b3)));
  assign y7 = (5'd10);
  assign y8 = ((p10<p13)?(!p6):(~&a2));
  assign y9 = (a3?b2:b2);
  assign y10 = (6'd2 * (a1&p2));
  assign y11 = {1{(~|({4{b0}}?{4{b2}}:((p6?a2:b1)<(a2?b2:b4))))}};
  assign y12 = {1{((((p14>=p11)>=$unsigned(p16)))==$signed(((b0<=p4)|(a3!==a3))))}};
  assign y13 = {1{{2{((a2==b3)&(p9&b0))}}}};
  assign y14 = (3'sd2);
  assign y15 = (((p1>>>p14)-(p10))+$unsigned((p10^p6)));
  assign y16 = (2'sd0);
  assign y17 = ((b2&a1)>>>$unsigned($signed(p8)));
endmodule
