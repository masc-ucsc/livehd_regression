module expression_00389(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(-2'sd0),(2'd2)};
  localparam [4:0] p1 = (^(((3'd2)?(3'sd2):(5'sd0))!=((4'd14)?(3'd2):(2'd3))));
  localparam [5:0] p2 = {{2{(-2'sd1)}},(~(4'd2))};
  localparam signed [3:0] p3 = {(&((((4'd3)>(3'd1))!==(~&((3'sd3)?(-5'sd11):(5'd15))))<<<({(5'sd1),(2'sd0)}?(6'd2 * (5'd13)):((3'sd2)<(-4'sd4)))))};
  localparam signed [4:0] p4 = ({1{(~^(-3'sd0))}}!==(!((|(2'sd1))>>>(4'd15))));
  localparam signed [5:0] p5 = {2{(-({3{(2'd0)}}&&((2'sd1)+(2'd1))))}};
  localparam [3:0] p6 = {{(4'd3),(3'd1),(-2'sd1)},(~^(3'd4))};
  localparam [4:0] p7 = ((-5'sd4)^(5'd29));
  localparam [5:0] p8 = (((3'd3)>>(4'd3))<<<((3'sd3)<(-2'sd1)));
  localparam signed [3:0] p9 = (({(4'sd5),(-4'sd1),(2'sd1)}>=(~|(2'sd0)))>(((2'sd1)<<(2'd0))&&((-5'sd5)?(2'sd0):(3'd4))));
  localparam signed [4:0] p10 = {3{(5'd30)}};
  localparam signed [5:0] p11 = ((3'd5)?(3'sd2):(4'd5));
  localparam [3:0] p12 = {(4'd1),(4'sd0)};
  localparam [4:0] p13 = (-((~&(~&(2'd0)))?((-2'sd1)?(-3'sd0):(5'd31)):(!(~&(3'sd2)))));
  localparam [5:0] p14 = ((~(((5'd10)!==(4'sd1))&((5'sd1)/(-4'sd6))))^((+(~&(|(5'd2))))^~(^(!((-5'sd14)>>>(3'd1))))));
  localparam signed [3:0] p15 = {{{{(2'sd1)}},{(4'd5),(3'd4),(2'd3)}},{{(3'sd3)},{(4'd12)},{(3'd3),(4'd13),(4'd2)}}};
  localparam signed [4:0] p16 = ((!(-(4'sd1)))+{4{(5'd16)}});
  localparam signed [5:0] p17 = {(5'sd11),(3'd6)};

  assign y0 = (($signed({p0}))?$signed((p1?p17:p1)):$signed({$signed(p14)}));
  assign y1 = (4'sd3);
  assign y2 = (~&(~^{(&{4{b5}}),(3'sd0),{1{(~^p8)}}}));
  assign y3 = ((b2>>b2)^~(a5>=b2));
  assign y4 = (|(b4));
  assign y5 = (5'd12);
  assign y6 = (~(+(~(~|(~(!((~&$signed(b4)))))))));
  assign y7 = (-((p2>>p10)==(!(p16>>p17))));
  assign y8 = (((5'd27)!=((5'd0)&(a0||a3)))+(-3'sd3));
  assign y9 = {{3{a4}}};
  assign y10 = ($unsigned(b1)|{4{a3}});
  assign y11 = {1{(({4{a1}}?(|p16):{p10})?((!p12)?{1{p5}}:(&p16)):{4{p0}})}};
  assign y12 = (~(p6!=b3));
  assign y13 = ((+(p11))^~$signed((&p14)));
  assign y14 = (((a4<<a4)>>(b4!==a4))!==((a1<<b3)|(a4^b0)));
  assign y15 = (((b5^~p13)?(b0>>>b4):{1{p14}})?{(p16?p13:p6),{p14},(^a5)}:(^(~(&$signed((p2<<p3))))));
  assign y16 = (~(((p9?b5:a2)?(p15?b1:b1):(~p17))?((a5-a1)===(a2>b3)):((~&(a1?a3:a4))!==(~&(b3?a5:a0)))));
  assign y17 = {((b5?a2:b2))};
endmodule
