module expression_00078(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd2)&(4'sd0))!=((2'sd0)&(5'sd0)))>(((5'd6)===(2'sd1))-{4{(5'd4)}}));
  localparam [4:0] p1 = (4'd12);
  localparam [5:0] p2 = ((-5'sd13)!=(5'd9));
  localparam signed [3:0] p3 = ({4{(3'd3)}}?((4'd0)?(2'd0):(-5'sd9)):((5'd17)?(5'sd4):(2'd1)));
  localparam signed [4:0] p4 = {{(-5'sd15),(3'd7),(5'd20)}};
  localparam signed [5:0] p5 = (((-2'sd1)==(3'sd2))>>((3'd0)?(2'd1):(4'sd7)));
  localparam [3:0] p6 = (-((~^(~((-3'sd1)||(4'd1))))!==(~(~^(&((2'd3)?(4'd0):(2'sd0)))))));
  localparam [4:0] p7 = {2{(~&{(5'd15),(-5'sd9)})}};
  localparam [5:0] p8 = {2{({(2'd3),(-4'sd7),(2'd2)}===(~|(5'sd2)))}};
  localparam signed [3:0] p9 = {(&{3{{(-4'sd1),(4'd7),(5'd9)}}})};
  localparam signed [4:0] p10 = {((-5'sd14)>>(5'd27)),((-3'sd3)&(5'sd4))};
  localparam signed [5:0] p11 = (&(3'sd1));
  localparam [3:0] p12 = ((~(^(-4'sd2)))===((2'd3)||(-3'sd1)));
  localparam [4:0] p13 = (((5'sd13)&(4'sd1))&((2'd1)>>(4'd9)));
  localparam [5:0] p14 = ((-3'sd2)!=(3'sd3));
  localparam signed [3:0] p15 = (3'd2);
  localparam signed [4:0] p16 = ({(5'sd15),(3'd7)}?((4'sd4)?(3'sd0):(3'd6)):(~^(4'd15)));
  localparam signed [5:0] p17 = {2{(6'd2 * (~(5'd4)))}};

  assign y0 = ((-{1{(~|((p11?p7:b1)-{1{b0}}))}})!={4{(&b3)}});
  assign y1 = (4'd4);
  assign y2 = ((&((b1-p11)==(b3<<<a2)))^((a1&&a4)%p10));
  assign y3 = {4{$unsigned($signed((a0^~a2)))}};
  assign y4 = (3'd3);
  assign y5 = ((5'd2 * $unsigned((~b1))));
  assign y6 = {4{(^p0)}};
  assign y7 = (4'd6);
  assign y8 = ((^(a4?a5:p17))<=(~(p7?p17:a5)));
  assign y9 = ({((p14?p0:b5)>>>$signed(p7))}>>>{{{p14}},(a5?p7:p7)});
  assign y10 = (~&(({1{p12}}?{1{p9}}:(p14>=p6))?((p5?p10:p8)|{3{p11}}):{4{(p12==p11)}}));
  assign y11 = {(5'sd14),(2'd3),(b4?b4:p15)};
  assign y12 = (3'd7);
  assign y13 = (5'd2);
  assign y14 = (|((^b2)?(a4?a5:p14):(2'd3)));
  assign y15 = {(p1||b3)};
  assign y16 = ((~&(p4&p16))?(p3?p11:p8):(p5?p1:p14));
  assign y17 = (($unsigned(a4)?(a2||a4):(a0===b3))?((a3?b2:a3)<<<(a0?p0:b3)):((b2||p12)>>>{4{a3}}));
endmodule
