module expression_00451(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(((-5'sd1)?(4'd9):(3'd0))?{1{((-3'sd0)?(2'd1):(3'sd1))}}:(((3'sd0)==(3'd2))===((-2'sd0)?(4'd10):(5'sd0))))}};
  localparam [4:0] p1 = ((|((3'sd1)?(-2'sd1):(3'sd3)))!=={(-3'sd3),(2'd0)});
  localparam [5:0] p2 = {{((6'd2 * (5'd8))>>>((3'sd3)||(3'sd3)))},(({(2'd3)}!=={2{(4'd14)}})==({(4'd8),(2'd3),(-4'sd0)}^{4{(4'd9)}}))};
  localparam signed [3:0] p3 = (-5'sd12);
  localparam signed [4:0] p4 = (5'd10);
  localparam signed [5:0] p5 = (((5'sd3)?(5'd15):(3'd2))*((2'd3)|(4'd15)));
  localparam [3:0] p6 = (((3'd3)?(4'd11):(3'sd1))===((-4'sd0)?(2'd2):(2'd0)));
  localparam [4:0] p7 = (-((~^(&(!{4{(4'd10)}})))&&((5'sd11)&&(!(4'sd7)))));
  localparam [5:0] p8 = {{(2'd1),{(3'd6),(-2'sd1),(-3'sd3)},{(4'sd2)}},(-5'sd12)};
  localparam signed [3:0] p9 = ((~|(5'd31))&&{(4'd11),(4'sd1)});
  localparam signed [4:0] p10 = (~(~&{(~&{(-(-5'sd15))}),(!{(4'd1),(3'd6)})}));
  localparam signed [5:0] p11 = (~^{(((4'sd7)!=(-4'sd3))>>{(2'sd0),(4'd10),(3'd1)}),(((3'd3)|(-5'sd5))^~(-(4'd1)))});
  localparam [3:0] p12 = {{{(~^(4'd12)),((4'd4)==(4'd7)),(~(5'd18))}},(~^(~^(+{((5'd25)==(2'd3))})))};
  localparam [4:0] p13 = {1{{({1{(4'sd0)}}?{(4'sd1),(3'sd0)}:{(-3'sd0),(2'sd0)}),{{{(4'd3),(3'd3)},{3{(-3'sd3)}}}}}}};
  localparam [5:0] p14 = (-4'sd2);
  localparam signed [3:0] p15 = (+{(-(!(-4'sd7))),((-2'sd0)?(5'd31):(5'd6)),((4'd4)?(5'd26):(-2'sd0))});
  localparam signed [4:0] p16 = (-(^(+(-(+((~|(~&(4'd12)))%(3'd6)))))));
  localparam signed [5:0] p17 = (!{{3{({(-4'sd5),(5'sd12),(3'd5)}&{(5'd29),(4'd12)})}}});

  assign y0 = (~^(|(((-(|p7))^(p9?b1:a3))?((+(p1?p6:p15))&(p8?p15:p2)):((|p15)?(b3?p13:a4):(p6?p1:a2)))));
  assign y1 = (((p4-p16)-(p9&&p5))&&((a3>=a5)!==(b1-a1)));
  assign y2 = {(5'd29),({p9}?{a2}:{p3}),($unsigned((p1>>>a0))^~(&(a1?p15:a0)))};
  assign y3 = (~^(^(|(|(5'sd11)))));
  assign y4 = (({1{b0}}?{1{p10}}:{b4})?{3{(3'd7)}}:{{4{{a1}}}});
  assign y5 = (-{2{(!b5)}});
  assign y6 = (~|(~(($unsigned((b5<=b3))!==(b2|b0))<=$signed(((!(!b0))+$signed((b5>>>b3)))))));
  assign y7 = $unsigned(((a3*b1)/a0));
  assign y8 = (({a1,a2}>>>{p3})-((p16==p8)!=(p14<<<b5)));
  assign y9 = (p3||b1);
  assign y10 = (|{((|(b1<<a4))==={a3,a3,a1})});
  assign y11 = (((5'sd7))>((~a0)^~(2'sd1)));
  assign y12 = (p1<=p17);
  assign y13 = {1{{4{{2{b1}}}}}};
  assign y14 = $signed((2'sd1));
  assign y15 = {2{(-4'sd6)}};
  assign y16 = {(4'sd3)};
  assign y17 = ((((p9||p11))^((a2>>>p17)>>(p5<<b5)))>>(($unsigned((p9^~p15))<=(4'd2 * p12))));
endmodule
