module expression_00328(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^{4{(&{1{(5'd7)}})}});
  localparam [4:0] p1 = (4'd12);
  localparam [5:0] p2 = (({3{(-2'sd1)}}-((2'sd0)>>>(-2'sd1)))-(((3'd0)<(2'sd0))>>>((-3'sd0)>>>(4'sd1))));
  localparam signed [3:0] p3 = ((-2'sd0)==((-5'sd9)!=(3'd7)));
  localparam signed [4:0] p4 = (3'sd1);
  localparam signed [5:0] p5 = (((~^{2{(-2'sd0)}})^{3{(4'd9)}})<<<({4{(4'd5)}}===(&((3'd1)>>>(-4'sd4)))));
  localparam [3:0] p6 = {({4{(3'sd0)}}>(!(2'd2))),{4{(2'sd0)}},((|(-5'sd13))?((2'sd1)?(-5'sd2):(4'd2)):((5'sd3)<<(4'd0)))};
  localparam [4:0] p7 = {((-4'sd7)&&(-2'sd0))};
  localparam [5:0] p8 = (({2{(3'd4)}}?(|(4'd9)):{3{(-3'sd1)}})&&(((2'd0)?(2'd2):(2'd0))?(&(2'd0)):{3{(3'd7)}}));
  localparam signed [3:0] p9 = (~&((^(~{1{(5'sd14)}}))&(-(|(~(2'd2))))));
  localparam signed [4:0] p10 = {3{{1{((4'sd7)<<<(2'sd1))}}}};
  localparam signed [5:0] p11 = ({(4'd15),(2'd2),(2'd2)}?((2'd1)?(-2'sd1):(-5'sd11)):((-2'sd1)?(-2'sd1):(5'd24)));
  localparam [3:0] p12 = (~|{{(-2'sd0),(4'd11),(2'd2)},{{(2'd3),(5'd30),(2'd3)}},(~&(~&(4'd13)))});
  localparam [4:0] p13 = (~(3'd2));
  localparam [5:0] p14 = (-(((2'd2)&&(2'd1))>=(!(~(2'sd0)))));
  localparam signed [3:0] p15 = {4{{1{((4'd13)+(3'sd1))}}}};
  localparam signed [4:0] p16 = (6'd2 * ((5'd27)|(4'd5)));
  localparam signed [5:0] p17 = {4{(!(-5'sd6))}};

  assign y0 = (~^((~^(|$unsigned(p11)))?((p0?p9:p0)):(p6?p6:p6)));
  assign y1 = ((p2?p16:p0)?{p5,p2,p9}:((p12&&p1)^(p12?p12:p8)));
  assign y2 = (((a3||p1)&(b2<b1))!={{p2,a3},(a4<<<p1)});
  assign y3 = $unsigned(((4'd1)&($signed((4'd7)))));
  assign y4 = $signed((5'd12));
  assign y5 = $unsigned($unsigned({2{({1{{4{p1}}}}<<((p8)||{1{p16}}))}}));
  assign y6 = ((a2!==a5)<<<{b1,a5});
  assign y7 = ((((-2'sd0)?(p16?p9:p13):(~p17)))<<<(4'd10));
  assign y8 = ((b5<a1)?(b3!==b3):(a1===b5));
  assign y9 = {3{$unsigned(b4)}};
  assign y10 = {1{{3{(a5>b2)}}}};
  assign y11 = (~&((5'd1)?(~|((&(p11?b5:p4))/a2)):(2'd1)));
  assign y12 = (~^$unsigned({3{({1{(p14>>>b3)}}-(b2+p6))}}));
  assign y13 = ((~|(5'sd15))?{(p4?p6:p3)}:(p8?b2:a5));
  assign y14 = (-(2'd0));
  assign y15 = (~&(~|((-p15)<<(a4+p13))));
  assign y16 = {2{(5'd16)}};
  assign y17 = {2{{2{p12}}}};
endmodule
