module expression_00570(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((((-4'sd5)?(5'sd2):(-4'sd6))>>((-3'sd2)?(2'd3):(4'd11)))^~(((4'sd2)&&(-4'sd3))^~((3'd3)?(5'd21):(3'd4))))&&({(-3'sd3),(4'sd1)}?(6'd2 * (3'd2)):((2'd1)+(5'd11))));
  localparam [4:0] p1 = ((4'd11)?(3'sd0):{1{((-4'sd3)!=(4'd13))}});
  localparam [5:0] p2 = (!((3'sd3)&{2{(2'd2)}}));
  localparam signed [3:0] p3 = ((((3'sd3)>>(-2'sd0))?(|(4'd13)):{2{(-5'sd3)}})!=({1{((2'sd1)?(4'sd1):(3'sd2))}}>=((-5'sd2)>>(3'sd3))));
  localparam signed [4:0] p4 = {1{(((4'sd3)?(2'sd1):(5'd22))?((2'sd0)?(4'd9):(-3'sd1)):((2'd1)+(4'd12)))}};
  localparam signed [5:0] p5 = (6'd2 * (4'd15));
  localparam [3:0] p6 = (5'd25);
  localparam [4:0] p7 = ((5'd15)>>(4'd1));
  localparam [5:0] p8 = (({(4'sd1),(5'd6),(3'sd0)}^~((3'd1)&&(2'd3)))||{{1{(4'sd2)}},(!(3'd6)),((3'd0)!==(3'd3))});
  localparam signed [3:0] p9 = (~&(~|(~^(&(~&(~|(^(-(+(3'sd2))))))))));
  localparam signed [4:0] p10 = (~|(|(5'd2 * ((4'd7)|(5'd12)))));
  localparam signed [5:0] p11 = (3'd5);
  localparam [3:0] p12 = (((2'd1)?(3'sd0):(2'd3))?(2'd2):{3{(4'd8)}});
  localparam [4:0] p13 = (|(~|(|((((2'd1)>(3'd7))&&((5'sd14)>(4'sd1)))?((-2'sd0)?(2'd0):(-4'sd1)):((~|(4'd9))>>((2'd0)-(5'd1)))))));
  localparam [5:0] p14 = (((((3'd0)?(2'd0):(2'sd1))===(~(-5'sd12)))>(-((4'sd5)!==(4'sd0))))==(!(((-2'sd0)+(-4'sd1))-(~&{(2'sd1),(3'd5)}))));
  localparam signed [3:0] p15 = ({3{((3'sd1)===(-4'sd6))}}^(-4'sd6));
  localparam signed [4:0] p16 = {{3{(4'sd6)}},((((4'd6)&(2'd2))>((5'd8)?(-4'sd6):(-4'sd1)))>={3{(3'd6)}})};
  localparam signed [5:0] p17 = ((3'sd0)%(4'd15));

  assign y0 = (-(({2{p16}}<=(^{p14,p4}))?((p16!=p7)?(p13<<p0):{p13,p3,p7}):(~|{(~|({4{p8}}+{3{p14}}))})));
  assign y1 = ((((a2===a5)<<<(b4?p12:a3))?$signed($unsigned({((b1&&a1))})):((a2>a4)?(a5||b4):{b4,p6})));
  assign y2 = (a1^b4);
  assign y3 = (({b2,b2}!==(b2^~a3))&{(a1<p6),(6'd2 * b2)});
  assign y4 = ({(~^b1),$signed(a2)}===(~(b1>>a4)));
  assign y5 = (((p13?p12:p10)-(p9&&p11))^{{p7,p1},$signed(p3),(p5^p14)});
  assign y6 = (((p15?p4:p6)?(~p6):(p17?p7:p13))?((p4>=a0)>>(p4?p9:p5)):(+((p11?p12:a5)&&(&(p8==p12)))));
  assign y7 = $unsigned((~&$signed((-4'sd7))));
  assign y8 = (!(4'sd7));
  assign y9 = ((((b1&a5)<(b5<b5)))===($signed(a1)?$signed(a3):(b2?a4:a3)));
  assign y10 = {p15,b3,b1};
  assign y11 = $unsigned(($signed((p11>p4))&$signed($signed(b0))));
  assign y12 = (4'd2 * (b2?p13:p13));
  assign y13 = (!((5'sd12)^~((-5'sd15)+(~^a1))));
  assign y14 = {2{p4}};
  assign y15 = (|(((~p8)?(p17?b4:p12):(~|a3))?(!(-(~|(~^(~p6))))):(&(~|(^(~(^a1)))))));
  assign y16 = (-5'sd4);
  assign y17 = (((p10>>>p13)>>>(a2))==({1{$unsigned($signed(b3))}}));
endmodule
