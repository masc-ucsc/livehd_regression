module expression_00593(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-2'sd1);
  localparam [4:0] p1 = ((2'sd1)<<<(-2'sd0));
  localparam [5:0] p2 = {((6'd2 * (~&(~&(3'd3))))&&(&(((3'd5)!=(-3'sd1))^((5'd13)+(2'sd1)))))};
  localparam signed [3:0] p3 = (!(|(~&{(!(-3'sd2)),(~&(4'd15)),{(2'd2),(-5'sd14)}})));
  localparam signed [4:0] p4 = (~&(4'd14));
  localparam signed [5:0] p5 = {4{(~^(!(-(4'd6))))}};
  localparam [3:0] p6 = (^{3{(~&(4'sd5))}});
  localparam [4:0] p7 = (+{(-5'sd9)});
  localparam [5:0] p8 = (((3'd0)!=(4'sd2))?((4'd6)^(2'sd1)):((3'sd0)^(4'sd2)));
  localparam signed [3:0] p9 = {(2'd3),(2'd0)};
  localparam signed [4:0] p10 = (^(5'd1));
  localparam signed [5:0] p11 = (4'd1);
  localparam [3:0] p12 = (|{{(|(5'sd6)),{(3'd2)},(2'd2)},{(+(5'd6)),((3'd0)?(4'd4):(-4'sd1)),(~^(2'd1))}});
  localparam [4:0] p13 = ((2'sd0)<<((5'd21)&&(-4'sd5)));
  localparam [5:0] p14 = (((4'd7)^(3'sd2))*((-5'sd14)&(5'd29)));
  localparam signed [3:0] p15 = (((-5'sd9)?(-3'sd0):(4'sd5))?{2{(3'd1)}}:{3{(5'd9)}});
  localparam signed [4:0] p16 = {3{{1{({1{(2'd1)}}=={1{(5'sd7)}})}}}};
  localparam signed [5:0] p17 = (((5'sd10)===(-3'sd0))?((-5'sd9)===(5'sd13)):(|(2'd2)));

  assign y0 = (((b5==b0))/b4);
  assign y1 = (~&(|{(({(a2^b3),(&a3)}==={(a3>b0),(b5>>b5)})>>((^{{p8,p3,p12}})<((a1<=b0)&&{a2,b3})))}));
  assign y2 = (p2&&p15);
  assign y3 = (((3'd3)!=(p14<b1))+(^((p0^~b5)&&(2'sd1))));
  assign y4 = ({b5,b4,a3}?(^(a1?b3:a2)):{b0,a2,b1});
  assign y5 = ((p8>=b5)?(+p16):{a1});
  assign y6 = $signed(((4'd2 * (b1?a2:a2))-((b1===b4)<(b5?p11:p3))));
  assign y7 = {4{((p0<=b0)>>{3{p9}})}};
  assign y8 = {4{(a3^~p10)}};
  assign y9 = (!(^(-(b4?a1:p11))));
  assign y10 = (!((~|(-(4'd2 * (-{p13}))))>>({p15,p2,a1}?(p10^p6):{(~|b0)})));
  assign y11 = (5'd21);
  assign y12 = {3{(p11?p4:p15)}};
  assign y13 = ((-5'sd13)^{3{{(4'd0)}}});
  assign y14 = ($signed((3'd7))>{($signed(a0)<{p6}),(~(p2>>>b2))});
  assign y15 = (((a1?p8:b3)&&(b5^~p2))<<<((~^b0)!=(p17?a5:p6)));
  assign y16 = (&({a5,p3,b5}?(a0?p8:a1):(a3?p7:a0)));
  assign y17 = $signed(a5);
endmodule
