module expression_00288(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'sd0)!=(-4'sd7))?((5'd30)<=(4'd2)):((-2'sd0)<<(2'sd0)))<(((5'd5)?(5'd4):(5'd13))?(5'd17):((2'sd1)?(5'd12):(-3'sd3))));
  localparam [4:0] p1 = {({2{{(3'd6)}}}&({4{(5'd12)}}==((-2'sd0)<=(5'd2))))};
  localparam [5:0] p2 = {4{{4{(5'd2)}}}};
  localparam signed [3:0] p3 = {4{{(4'd0),(5'd0),(5'd0)}}};
  localparam signed [4:0] p4 = {((2'd1)<(2'd3)),{(5'd7),(-3'sd3)}};
  localparam signed [5:0] p5 = ((((5'd8)-(-2'sd1))&((5'd21)<<<(3'd1)))>>(((-3'sd1)>>>(3'sd0))!==((4'd8)?(-5'sd2):(5'd6))));
  localparam [3:0] p6 = {2{(2'sd0)}};
  localparam [4:0] p7 = ((-3'sd3)?(~^(-2'sd1)):(~^(5'sd6)));
  localparam [5:0] p8 = ((4'd8)?(5'sd6):(3'd6));
  localparam signed [3:0] p9 = {((5'd20)&&(2'sd1)),{(5'sd14)}};
  localparam signed [4:0] p10 = (((5'sd13)?(3'sd1):(-3'sd2))^~{((4'd9)?(4'd6):(4'd6)),{(3'd2),(-3'sd0)}});
  localparam signed [5:0] p11 = (((4'sd0)<<<(3'd5))!=((5'sd13)*(2'sd1)));
  localparam [3:0] p12 = (((-3'sd3)<<((3'd0)?(-4'sd0):(5'd0)))?(((5'sd0)?(2'd0):(4'sd3))&&((5'd14)%(-4'sd6))):((2'sd1)?(5'd27):(3'd3)));
  localparam [4:0] p13 = {1{({((4'd10)?(5'd13):(2'sd0))}||{2{{4{(3'd2)}}}})}};
  localparam [5:0] p14 = ({2{((3'd1)>(3'd0))}}-{4{((3'd3)!=(-2'sd0))}});
  localparam signed [3:0] p15 = (((4'd2)+(5'd23))^~{3{(-2'sd0)}});
  localparam signed [4:0] p16 = (4'd15);
  localparam signed [5:0] p17 = ((3'd3)!==(-5'sd0));

  assign y0 = $unsigned({3{($unsigned((a1&p16)))}});
  assign y1 = $signed((((4'd2 * p12)<<<$signed(p16))<=(|(3'sd3))));
  assign y2 = (4'sd1);
  assign y3 = ((p13?a3:p8));
  assign y4 = (((((b0>b5)*(b3<<<b1))))|$unsigned((($unsigned(a3)&&(b4))>((b1)^$unsigned(p10)))));
  assign y5 = $unsigned((6'd2 * a0));
  assign y6 = ({1{(((5'sd3)>={2{a4}})!==$unsigned((a2-b1)))}}||(-3'sd1));
  assign y7 = {2{{1{{1{{1{{4{p13}}}}}}}}}};
  assign y8 = ((a1?a0:a0)|{{3{b5}},(a1)});
  assign y9 = {2{$unsigned(({2{a0}}?$unsigned($unsigned(p10)):(p7?b4:a2)))}};
  assign y10 = {((4'sd2)<<(5'd29))};
  assign y11 = ((b2?a0:p6)?(a4?a0:a1):(b3?b4:b0));
  assign y12 = (-2'sd1);
  assign y13 = (+({{$unsigned((2'sd1)),(a4>=b5),{(b2<b4)}}}===(+{3{(2'd1)}})));
  assign y14 = (~&(((-3'sd1)<<<(-3'sd3))>>>(4'sd2)));
  assign y15 = (~&(~|(~(+(|(&a2))))));
  assign y16 = ((a4^~b0)<{3{b4}});
  assign y17 = ($unsigned(((p8<=p14)<(-5'sd11)))^~{(p9>=p2),{p16,p1},(p4<p1)});
endmodule
