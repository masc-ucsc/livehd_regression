module expression_00601(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{4{((-5'sd5)>>(5'd27))}}};
  localparam [4:0] p1 = {{{(-2'sd0)},{(3'd6),(3'd3),(4'sd0)},{(4'd13),(3'd5),(3'd6)}},(+(((-4'sd1)<=(3'sd3))!==(-2'sd0)))};
  localparam [5:0] p2 = (-((-4'sd0)<<<(-2'sd0)));
  localparam signed [3:0] p3 = (^((2'd2)>(-4'sd6)));
  localparam signed [4:0] p4 = (+((((5'sd14)>=(5'sd13))^((2'd0)<<<(3'd0)))^~(((3'sd0)===(2'd1))||((4'sd7)&&(4'sd5)))));
  localparam signed [5:0] p5 = (2'd1);
  localparam [3:0] p6 = {(~&((3'd5)?(2'd0):(5'sd13))),((3'd2)?(3'sd2):(3'sd3)),(~((4'd11)?(5'd26):(3'sd1)))};
  localparam [4:0] p7 = {4{(-2'sd0)}};
  localparam [5:0] p8 = {2{{2{(-3'sd2)}}}};
  localparam signed [3:0] p9 = (-2'sd0);
  localparam signed [4:0] p10 = {{{{(-4'sd4)},((3'd3)<<<(5'd14))}},{{2{{4{(-3'sd0)}}}}},{4{(5'd0)}}};
  localparam signed [5:0] p11 = ((3'd3)|(4'd8));
  localparam [3:0] p12 = ((~(~&((-(2'd1))>>>((4'sd3)>=(5'sd11)))))>((~&(&(-5'sd7)))||((4'd3)/(-2'sd0))));
  localparam [4:0] p13 = (({(-5'sd9),(2'd1)}|(~(2'sd1)))!=={(^(!(3'sd1)))});
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = (~|({4{((3'sd1)?(2'd1):(2'd1))}}<={2{((-2'sd1)==(4'sd5))}}));
  localparam signed [4:0] p16 = (5'd2 * ((3'd0)===(2'd2)));
  localparam signed [5:0] p17 = ({4{(5'd17)}}^~{2{((4'sd2)?(3'd2):(5'd2))}});

  assign y0 = {2{a2}};
  assign y1 = ((~&((p8?b2:b0)?(p12?b2:b0):(&b3)))>=(!(~(|(+(a0?p2:a0))))));
  assign y2 = ({((p9<<b5)||{3{a4}}),{p14,a1,a1}}<({{4{b0}},{4{b2}}}==((b5+b3)>>(6'd2 * b2))));
  assign y3 = ({3{a5}}<<((^(a5>>b5))));
  assign y4 = {4{{1{b1}}}};
  assign y5 = ((-(~|{(~a4),(|b3)}))!=={{((a3!==a4)^(a3<<<a5))}});
  assign y6 = {3{{2{p0}}}};
  assign y7 = (^(((a4>=a0)<<<(|a2))?(-(|(p15>>>b4))):((-a1)+(b3>>b3))));
  assign y8 = {(-(a3?b3:b0))};
  assign y9 = ({b2,p9,a0}-(~&{a0,b3}));
  assign y10 = {2{{{2{a4}}}}};
  assign y11 = ({2{a4}}?{1{a4}}:{2{b2}});
  assign y12 = (^({2{(&(p2?a3:p10))}}^~(~^({1{(~|p8)}}>>(p10<<p10)))));
  assign y13 = ((!((!(p6+b0))|((p14-p16)|(~&p13))))>(-{4{{1{a0}}}}));
  assign y14 = (b5^p4);
  assign y15 = (((b1<=a0)%p0));
  assign y16 = $unsigned(b5);
  assign y17 = (p6+p7);
endmodule
