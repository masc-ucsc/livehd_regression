module expression_00309(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{(((2'd0)<<(2'sd1))&&((-5'sd1)&(5'd17)))}};
  localparam [4:0] p1 = {2{(((3'd4)==(3'd0))|(-(4'd3)))}};
  localparam [5:0] p2 = {1{(((3'sd0)!==(3'd7))!==((4'd8)!=(-3'sd1)))}};
  localparam signed [3:0] p3 = (3'd1);
  localparam signed [4:0] p4 = ((5'd19)||(-3'sd3));
  localparam signed [5:0] p5 = {(|{(-5'sd7),(2'd3)}),(~^{(5'd10),(5'sd14)}),{(~^(5'd28))}};
  localparam [3:0] p6 = ({3{(-2'sd1)}}?((-3'sd1)?(2'd2):(5'd11)):((2'sd1)===(4'd12)));
  localparam [4:0] p7 = (~((5'd16)>=(~(&(3'd1)))));
  localparam [5:0] p8 = (((&(~^(5'd20)))&&(~&((-5'sd3)|(5'sd7))))-(((5'd6)<=(2'sd0))>>>(-((2'sd0)<<<(5'sd3)))));
  localparam signed [3:0] p9 = (((|(~|(2'd3)))>>((5'sd8)^(-3'sd0)))!=={{(-5'sd9),(-3'sd3),(4'sd6)},{1{{(4'sd0)}}}});
  localparam signed [4:0] p10 = ((4'sd2)>=(4'd13));
  localparam signed [5:0] p11 = (((3'd1)?(5'sd0):(4'd1))/(5'sd0));
  localparam [3:0] p12 = {(((5'd0)===(5'd19))<<<((-3'sd1)+(5'd5)))};
  localparam [4:0] p13 = (2'd3);
  localparam [5:0] p14 = (~&{(((~&((-4'sd0)!==(2'sd0)))===(~&{(-3'sd3)}))<=(!(((5'sd6)!=(5'sd9))!={(4'd12),(2'd1),(5'd25)})))});
  localparam signed [3:0] p15 = (|(((3'd3)<<<(3'd1))<=(-((3'd1)>(4'd11)))));
  localparam signed [4:0] p16 = (5'd2 * {(~^(5'd28))});
  localparam signed [5:0] p17 = (-({((2'd1)?(-2'sd0):(5'sd3)),(!(-3'sd1)),((4'd12)?(-5'sd13):(-5'sd5))}>=((|(3'd3))?((5'd13)>>>(5'd15)):((3'd6)>(4'd15)))));

  assign y0 = (p7?p12:p5);
  assign y1 = {{a2,p2,a0},((p8)|{a1,p15}),({a3,p17}==(p8^~p9))};
  assign y2 = (2'd2);
  assign y3 = ((({3{b4}}==(~^b3))!=(|{3{b1}}))==({1{$unsigned((^a5))}}!==$signed({(b2^~a5)})));
  assign y4 = ($signed((b0/b0))?(a0?a0:b2):$unsigned((b2<a2)));
  assign y5 = (2'd2);
  assign y6 = ((-2'sd1)^~(+p6));
  assign y7 = ((p7-b2)>{3{b5}});
  assign y8 = ((-3'sd2)?(b2?p6:b3):(-5'sd4));
  assign y9 = (p5);
  assign y10 = ((((5'd2 * a1)>>(-5'sd4))<=((p16|b0)+(-3'sd3)))<(5'd2 * (p8>p14)));
  assign y11 = {{p16,p11},(!(5'd2 * b2))};
  assign y12 = {4{{2{(a0&&b3)}}}};
  assign y13 = (((4'd11)<<{a3,p8,p0})|{a0,b1,p0});
  assign y14 = {2{((+a4)?(~&p11):(~^p16))}};
  assign y15 = (6'd2 * b1);
  assign y16 = (a0?p8:b3);
  assign y17 = ({2{({4{b4}}|(a1>=p13))}}>>>((p4>>>p1)?{2{b5}}:(p1<=a3)));
endmodule
