module expression_00561(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{1{{2{{2{(4'sd0)}}}}}}}};
  localparam [4:0] p1 = (4'sd4);
  localparam [5:0] p2 = {(-(+(5'd26))),{(-3'sd3),(5'd17)},(&{2{(4'd5)}})};
  localparam signed [3:0] p3 = ((((5'd22)^~(-3'sd2))<<(^((2'd2)+(5'd16))))==={4{(~|(5'd4))}});
  localparam signed [4:0] p4 = (!(((3'd1)&&(4'sd3))>>{2{(-2'sd1)}}));
  localparam signed [5:0] p5 = (5'd18);
  localparam [3:0] p6 = (4'sd2);
  localparam [4:0] p7 = (((5'd27)<=(-3'sd3))*(~^((3'd7)*(-5'sd2))));
  localparam [5:0] p8 = ((((2'd0)||(4'd11))?((5'd31)==(4'sd3)):{(5'd8),(-4'sd0),(4'd11)})||(((2'sd0)>>(-5'sd6))>=((-5'sd2)>>>(3'd0))));
  localparam signed [3:0] p9 = ((-5'sd8)<<((5'd13)?(-2'sd1):(2'd3)));
  localparam signed [4:0] p10 = {(5'd2 * (~(6'd2 * (3'd2))))};
  localparam signed [5:0] p11 = ((((3'd1)<=(3'sd1))||((2'sd0)<=(5'd12)))<<<(((4'd5)|(3'sd0))!==((-2'sd0)|(4'sd3))));
  localparam [3:0] p12 = ((~&{(-3'sd2),(5'd19)})>(|{{(2'd2),(-4'sd4),(5'd10)}}));
  localparam [4:0] p13 = ((~&({(4'd4),(5'd12),(4'sd4)}>=(-(3'sd3))))?({(2'sd0)}&&(-3'sd0)):(((4'd12)?(4'd15):(-3'sd0))&&(^(4'd1))));
  localparam [5:0] p14 = ((4'd10)^~(2'd2));
  localparam signed [3:0] p15 = {2{{3{(-3'sd1)}}}};
  localparam signed [4:0] p16 = (~((5'd26)^~(5'sd2)));
  localparam signed [5:0] p17 = ((3'd3)-(3'd1));

  assign y0 = (2'd2);
  assign y1 = (|((-(~((~p12)|(~a3))))?(!(+(~|(a1?b4:a0)))):(~^((^b5)!=(p4?b3:p14)))));
  assign y2 = {1{{1{(b5&&p13)}}}};
  assign y3 = (+{3{$unsigned(({p1,a1}!=(b1)))}});
  assign y4 = $unsigned($signed((+p2)));
  assign y5 = {2{(-4'sd2)}};
  assign y6 = ({{a4,a2,a0},{p17,p10},(a5==a0)}>(~^(+{(~|((-b2)>>(a4||p15)))})));
  assign y7 = (((-4'sd6)||(~(a3?a1:p14))));
  assign y8 = ((p14>>p17)>{4{b1}});
  assign y9 = (~(2'sd1));
  assign y10 = (+(~({p13,p3,p1}?{1{{{p3}}}}:{4{p3}})));
  assign y11 = {4{{p4,b1,p16}}};
  assign y12 = ((+((p10>p3)+(~|b4)))?(-((a5===a1)!=(p14?p3:p17))):((p17?p8:p15)?(|b1):(~^p5)));
  assign y13 = (~(5'd28));
  assign y14 = {2{({b2,b1,a4}>=(5'd2 * b2))}};
  assign y15 = (5'd27);
  assign y16 = (((b2?a0:a2)!=((p9<b5)==(a2-b5)))<((p15!=b4)?(a2!==b5):(a4&&b4)));
  assign y17 = ((p15<<p12)<<(p5?p15:p7));
endmodule
