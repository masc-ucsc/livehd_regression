module expression_00216(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(~^(+(^(!(-(|(~&(&(5'd22))))))))));
  localparam [4:0] p1 = ((((-3'sd3)?(2'd0):(3'sd1))/(3'd2))?((~|(-4'sd2))&((-2'sd0)>=(3'sd0))):(~((5'd4)?(2'd0):(2'd3))));
  localparam [5:0] p2 = (-(~(~^(~((-(((5'd16)>>(-2'sd1))||((2'sd1)<=(5'sd0))))>>>(~^((~|(5'sd15))<(|(2'd0)))))))));
  localparam signed [3:0] p3 = ((4'sd5)?(-5'sd11):(2'sd0));
  localparam signed [4:0] p4 = (5'd12);
  localparam signed [5:0] p5 = ((-4'sd1)?(2'd2):(2'sd1));
  localparam [3:0] p6 = (((~&(~^(3'd7)))?((3'd3)?(-3'sd0):(4'd14)):(~|(+(5'd27))))^(!(&((~^(-(2'd2)))===((4'd5)>=(4'd11))))));
  localparam [4:0] p7 = (&(-5'sd2));
  localparam [5:0] p8 = (!(5'sd4));
  localparam signed [3:0] p9 = {1{({1{{1{((3'd7)<<<(3'sd0))}}}}!=(-3'sd3))}};
  localparam signed [4:0] p10 = {3{(-3'sd1)}};
  localparam signed [5:0] p11 = (-(2'd1));
  localparam [3:0] p12 = (~(~^(!(~^(|(~|(^(^(|(^(!(&(|(!(~(4'd3))))))))))))))));
  localparam [4:0] p13 = (+(+(-{(-{(&(3'd4)),{(3'd0)},(|(-4'sd7))})})));
  localparam [5:0] p14 = ({1{({1{(-2'sd1)}}<<((2'd0)!==(4'd8)))}}^~({2{(5'd14)}}^{3{(2'sd1)}}));
  localparam signed [3:0] p15 = ((4'd0)<(4'sd2));
  localparam signed [4:0] p16 = (!((((-3'sd1)*(5'd9))||((-2'sd1)?(3'd6):(5'd0)))<<<(((5'd8)^~(-5'sd2))?(!(4'd4)):((-4'sd5)!=(4'sd0)))));
  localparam signed [5:0] p17 = (^(~&(5'd2 * (4'd5))));

  assign y0 = {4{((a2&&p3)>=(4'd2 * p2))}};
  assign y1 = (~(p11-p11));
  assign y2 = {2{p2}};
  assign y3 = (($signed(a1)?(~&a3):(p3?a0:b4))>>>$unsigned($signed(((~^b4)+(p15?a1:a4)))));
  assign y4 = ({4{(a0!=p3)}}!={2{({2{b4}}>(6'd2 * a2))}});
  assign y5 = ({3{(a2>>b5)}}===((b1===a3)>=(a1<<a5)));
  assign y6 = ($signed($signed((~|((p16>>>p6)!=(p12-p9)))))+$signed((~(~|((p16>>p7)>>>(p13-p9))))));
  assign y7 = ({(-5'sd5),$signed({p6,p9}),{1{(p14&p15)}}}>=(-2'sd1));
  assign y8 = $unsigned((($unsigned((^(p7||p11)))|((!p7)!=(p6<<<p13)))));
  assign y9 = (2'd2);
  assign y10 = (b3?a2:b2);
  assign y11 = {4{(~^(p0>>b1))}};
  assign y12 = $unsigned(($signed(($unsigned((b2?a5:b3))?((b0?b0:a3)?(b2-a4):{2{a1}}):{3{(p9?b5:b5)}}))));
  assign y13 = $unsigned({a4,b5,a5});
  assign y14 = (~|(((5'd22)|((~^b1)<<(&p17)))));
  assign y15 = (((p13+p9)>(-3'sd3))^~(4'd6));
  assign y16 = $signed($signed($signed((($signed({3{p10}}))?(-({3{p12}}?(p3?p6:p6):{4{p3}})):{4{{2{p13}}}}))));
  assign y17 = $unsigned($signed(({{$signed((a4<a0)),{(b0>a0)},(a4||b3)}}||(({({b0,a4})}||((4'd2 * a0)>>{b1,b3,a4}))))));
endmodule
