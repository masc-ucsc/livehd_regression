module expression_00206(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-4'sd0)&(-2'sd1));
  localparam [4:0] p1 = ((+(^(3'd5)))&&(^{1{(5'sd4)}}));
  localparam [5:0] p2 = (~^(6'd2 * ((2'd0)^~(5'd24))));
  localparam signed [3:0] p3 = ((-3'sd2)=={4{(-5'sd3)}});
  localparam signed [4:0] p4 = ((((5'd6)<=(3'sd3))<<<{(2'd0),(4'sd4)})<<{((5'd6)<<<(-2'sd1)),{(-2'sd1)},{(-5'sd0)}});
  localparam signed [5:0] p5 = ({(~&(-2'sd1)),((3'd3)<<(4'd15)),{(2'd1),(3'd4)}}^(+{{(3'sd3),(3'd2)},((2'd3)!==(-4'sd4))}));
  localparam [3:0] p6 = ((3'd4)?(5'd30):(2'sd0));
  localparam [4:0] p7 = (2'd2);
  localparam [5:0] p8 = {4{(2'd3)}};
  localparam signed [3:0] p9 = (-3'sd2);
  localparam signed [4:0] p10 = (5'd2 * (4'd13));
  localparam signed [5:0] p11 = {((3'sd2)<<<(2'sd0))};
  localparam [3:0] p12 = ((!(5'sd2))>=((2'sd1)<(3'd4)));
  localparam [4:0] p13 = {4{{2{{(2'd0),(-2'sd1)}}}}};
  localparam [5:0] p14 = (+((-3'sd0)&(5'd17)));
  localparam signed [3:0] p15 = {1{(((-3'sd1)?((5'd5)<(2'd2)):((2'd1)>>>(3'sd3)))<{3{{4{(4'd2)}}}})}};
  localparam signed [4:0] p16 = (((6'd2 * (3'd1))>(!(5'd2 * (3'd0))))>>{(~&(4'd13)),((4'd0)==(3'sd1)),((2'd1)>=(2'sd0))});
  localparam signed [5:0] p17 = (~&((-4'sd0)!==(2'sd0)));

  assign y0 = {{4{{3{p17}}}}};
  assign y1 = ((((p10>>>p1))?(p12|p11):(p14?p1:p10))&(((p5<p10)^~(p12-p16))>>(a4?p13:p12)));
  assign y2 = (|((-(4'd8))&(5'd5)));
  assign y3 = (5'd16);
  assign y4 = (((p10<<p12)>=(p17+p13))!=((p6?p4:p12)>>>(+(b0?p16:p6))));
  assign y5 = (((~^$signed(b4))==$signed((+a1)))?((b3&&b5)===(b1>>b1)):((a1?a1:a5)?(p15+a4):(b2?b0:b1)));
  assign y6 = (5'sd7);
  assign y7 = (-2'sd0);
  assign y8 = (&(!{(+p17),{p7,p16,p10},(&p11)}));
  assign y9 = (($signed((p5<p9))=={3{p1}})>$unsigned(($signed((~(3'd4)))>(3'd0))));
  assign y10 = (!(4'd2 * {4{p14}}));
  assign y11 = (5'd29);
  assign y12 = (({(b4>=b0)}?$signed((a0!=b4)):(a2!==a5))!==({(a0?a2:a5),(4'd2 * b2),(b2<<<a2)}^~((a2?a1:a5)>=(a1?a5:a0))));
  assign y13 = {(4'd2 * {a2,a0}),{3{{2{b2}}}}};
  assign y14 = ((~&(a2?b2:b5))|(4'd2 * b0));
  assign y15 = (5'd2 * {a2,b2,b0});
  assign y16 = (({3{p9}}<<<(+a4))?((p2||p5)^~(~&p8)):(p5?p14:p10));
  assign y17 = (2'sd0);
endmodule
