module expression_00478(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd0)^~(-5'sd13))&((4'sd3)<<(4'd13)));
  localparam [4:0] p1 = {4{(5'd12)}};
  localparam [5:0] p2 = ((((-5'sd3)<<<(2'd1))^((-5'sd14)<<<(4'd10)))-(((-2'sd0)^~(-4'sd7))|(~(5'd3))));
  localparam signed [3:0] p3 = (&(+(|(5'd13))));
  localparam signed [4:0] p4 = (~^{3{(!(5'sd2))}});
  localparam signed [5:0] p5 = (~^({((-5'sd10)^(-3'sd2)),((-2'sd0)<<<(5'd25))}+{{(-3'sd0),(2'd1)},((-2'sd0)<=(5'd30)),(-(5'd14))}));
  localparam [3:0] p6 = (((4'd4)?(-4'sd3):(4'd10))?((-2'sd0)?(-2'sd1):(5'sd0)):((-4'sd6)?(3'd6):(-2'sd0)));
  localparam [4:0] p7 = {({2{(-2'sd0)}}||{((5'sd3)&&(3'd4))}),{((3'd7)^~(-5'sd6)),(-5'sd15),((-3'sd2)<=(2'd2))}};
  localparam [5:0] p8 = (-3'sd1);
  localparam signed [3:0] p9 = (-(-2'sd1));
  localparam signed [4:0] p10 = {2{((-3'sd0)+(5'd31))}};
  localparam signed [5:0] p11 = ((~|((5'sd12)?(4'sd5):(4'sd5)))^(+(~&(4'sd6))));
  localparam [3:0] p12 = {2{(-4'sd3)}};
  localparam [4:0] p13 = (((^(3'd4))?((4'd2)?(2'sd0):(-4'sd6)):((-2'sd0)?(-3'sd3):(4'd0)))?(~&(-(+((4'd12)&(5'sd9))))):(~^(((3'sd1)?(3'd7):(5'sd6))+((4'd12)+(-2'sd0)))));
  localparam [5:0] p14 = {3{(~^(5'sd8))}};
  localparam signed [3:0] p15 = {{(-5'sd9),(3'd1),(3'sd2)},{(-4'sd6),(2'd2),(-5'sd6)},{(4'd7),(-2'sd0),(5'd30)}};
  localparam signed [4:0] p16 = (((-4'sd7)^(4'sd0))>>((-5'sd10)<<<(2'd3)));
  localparam signed [5:0] p17 = (~^(((~|(4'd8))<=(-(3'd4)))<((~&(2'd2))!=(~&(-3'sd0)))));

  assign y0 = $unsigned($unsigned((((($signed({a0,p13,a5}))=={b1,p10,a5})>>>$unsigned($unsigned($signed({(p13>=p11),$unsigned((a4))})))))));
  assign y1 = (^(!(~&(!$signed({(((~p12)?(^p7):(p8))),{{(b0?a0:p17),{b2,p17}}}})))));
  assign y2 = ((!(-5'sd5))==={1{((({a0,b3}^~$unsigned(b5))!==(5'd2 * $unsigned(b1))))}});
  assign y3 = (((+((5'sd3)<=(b3==b5)))&((5'd2 * a2)^(4'sd2)))===(-4'sd6));
  assign y4 = (b1<=b4);
  assign y5 = {(~{(~&p8),{3{a5}},{1{p7}}})};
  assign y6 = ((((p14>p0)>>(p10==p10))||(~|$unsigned((p11^p2))))|((p13<=p15)%p5));
  assign y7 = $unsigned(((p7?p12:p12)?{a4,a1}:$signed(a0)));
  assign y8 = {p11,p16,b0};
  assign y9 = (!(!((^$unsigned((!(^$signed((p15||p16))))))|((~|(^p8))>>$signed((~&p7))))));
  assign y10 = (({a0,b4}>={b4,a3})^((b0|b4)^(4'd2 * b1)));
  assign y11 = (a4!==b5);
  assign y12 = {1{(-(~^((p2)?(p1):(p1))))}};
  assign y13 = $unsigned(({b4,b3,a2}?(a0?b4:b2):(p3>>>p0)));
  assign y14 = {({a1}?{a2}:(5'd2 * b1)),(+{2{(b5<=b3)}}),(+((-p2)^(a4^p8)))};
  assign y15 = {3{{1{(~&(-(!p7)))}}}};
  assign y16 = {$unsigned(a1),(-4'sd5),(p6)};
  assign y17 = ((-3'sd3)?{{p2,p4},{{p17,a0}}}:((b3?p11:b4)?(b4?p12:p12):(b1!==a3)));
endmodule
