module expression_00692(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(~|(^(-2'sd0))));
  localparam [4:0] p1 = {((-2'sd0)^(4'd3)),((5'sd5)&(5'sd7))};
  localparam [5:0] p2 = (({(3'd7)}^((3'd1)-(4'd11)))&{3{(-2'sd1)}});
  localparam signed [3:0] p3 = (4'd2 * (~((3'd7)>>>(5'd17))));
  localparam signed [4:0] p4 = (|{(5'sd13),(3'd4),(4'sd3)});
  localparam signed [5:0] p5 = ((4'd8)-(((2'd1)!=(3'sd3))&&(3'd6)));
  localparam [3:0] p6 = (((-2'sd1)?(5'sd9):(2'd1))*((-3'sd2)?(2'sd1):(5'd30)));
  localparam [4:0] p7 = (-5'sd10);
  localparam [5:0] p8 = (^{(!((4'sd1)^~(2'd1))),((5'd20)>>(-5'sd3)),{(3'sd1),(-5'sd12)}});
  localparam signed [3:0] p9 = (((&(4'sd4))<=(3'sd0))<=(2'd0));
  localparam signed [4:0] p10 = (5'd9);
  localparam signed [5:0] p11 = (&((-2'sd1)?(2'd0):(5'd25)));
  localparam [3:0] p12 = (|(!({{(3'sd2)},{(-5'sd13),(-4'sd5),(5'd13)}}>>(5'd2 * {(2'd1),(4'd15)}))));
  localparam [4:0] p13 = ((((5'd11)|(-4'sd1))?((5'sd8)>(-4'sd0)):((2'd2)?(2'd1):(-5'sd5)))!={(~&(-2'sd0)),(^(-3'sd1)),(~^(3'd2))});
  localparam [5:0] p14 = (&(5'd4));
  localparam signed [3:0] p15 = ((4'd8)?((|(2'sd0))?((-3'sd1)?(3'sd3):(3'd5)):(5'd21)):(((5'sd15)?(4'd9):(3'd0))<=((2'd0)?(4'd11):(-4'sd7))));
  localparam signed [4:0] p16 = (((3'd6)<(2'sd1))?(2'd0):((2'sd0)?(4'd8):(5'sd0)));
  localparam signed [5:0] p17 = ((3'sd0)&&(3'd0));

  assign y0 = (((a2>b2)!=(a0^a0))>((a1||a4)>(a5*b4)));
  assign y1 = ({a0,b0}!=(4'd2 * b2));
  assign y2 = ((&{2{(4'd3)}})>((6'd2 * b0)||(a4&&p9)));
  assign y3 = (({2{a4}}^{1{a0}})>>>{{a3,p9,b5}});
  assign y4 = {((((b1?b0:p7)<<<(p11!=p12))))};
  assign y5 = (((!(b4===b2))>>>$signed({3{p14}}))>=$unsigned($signed((-(|(a4!==b1))))));
  assign y6 = ((~|a2)!==(b3||b3));
  assign y7 = (5'd4);
  assign y8 = ((5'sd3)==(~^((a3!==a1)?(p4?p3:b1):(!p4))));
  assign y9 = ({(-((+p14)>>>(p2&p3))),{1{{2{(4'd2 * p7)}}}}}^({((&p7)<={1{p8}}),(~(p11&p6))}));
  assign y10 = (((^(+b5))-(b4?b2:b4))&((~|(~($signed(p7)<(b0||p17))))));
  assign y11 = ((((-5'sd1)+{b3,b1,p0})<<(~&(4'd2 * b0)))>>>(-((b3>>>b0)>{a3,p0})));
  assign y12 = {3{{1{a2}}}};
  assign y13 = {(p2<<p4),(p16==p5),(&(p2&&p5))};
  assign y14 = (^(|$unsigned((4'd0))));
  assign y15 = {(((a2&a3)?{b3,p5,b5}:(p12?b2:a2))>({p14,b5}?{b0,a5}:(b2?p5:p5)))};
  assign y16 = ((p4<<<p3)&&(p16^p2));
  assign y17 = (2'd2);
endmodule
