module expression_00592(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(4'sd1)}};
  localparam [4:0] p1 = {1{{3{(2'd2)}}}};
  localparam [5:0] p2 = (-2'sd1);
  localparam signed [3:0] p3 = (((-2'sd0)?(4'd8):(-5'sd13))?(&(3'd7)):((5'd22)?(3'd1):(3'sd0)));
  localparam signed [4:0] p4 = (((-4'sd5)?(-5'sd7):(-2'sd1))?(4'd2 * (3'd2)):(6'd2 * (5'd0)));
  localparam signed [5:0] p5 = (((4'sd6)?(4'sd3):(4'd13))?{1{(~^((3'd5)?(-2'sd0):(2'd3)))}}:(-(-((5'sd14)?(-4'sd5):(3'd4)))));
  localparam [3:0] p6 = ({{(4'd11),(3'd7),(4'd9)},(-(3'd1)),((-5'sd3)?(5'sd8):(2'd3))}?(^((5'd11)?(3'd5):(3'd6))):{4{(2'd1)}});
  localparam [4:0] p7 = ({4{(4'd7)}}&{(3'd5),(4'sd7),(5'd28)});
  localparam [5:0] p8 = {((-5'sd5)?(-(-4'sd7)):{(-4'sd6),(5'sd7)})};
  localparam signed [3:0] p9 = (4'd2);
  localparam signed [4:0] p10 = (2'sd1);
  localparam signed [5:0] p11 = (2'd3);
  localparam [3:0] p12 = (~^(&((5'd30)==(3'd1))));
  localparam [4:0] p13 = (((2'd0)<<(-2'sd0))=={(3'd5),(-3'sd3)});
  localparam [5:0] p14 = (-(5'd12));
  localparam signed [3:0] p15 = ({1{{3{((2'd3)^(3'sd2))}}}}>={1{({{(5'sd14),(2'd1),(2'd1)}}|{4{(-4'sd2)}})}});
  localparam signed [4:0] p16 = (3'sd2);
  localparam signed [5:0] p17 = (2'd1);

  assign y0 = ((~&((~&b0)===(b5&&b1)))?((b1?a1:a2)?(b1&&a3):(^a5)):((&a0)<<<(a3?p6:b1)));
  assign y1 = ({p7}|(~|a0));
  assign y2 = {2{{3{$signed(a4)}}}};
  assign y3 = ((a3<=b0));
  assign y4 = ((|{1{{(&$unsigned({3{p0}}))}}})^~$signed({1{({p8,p15}||(a0^~a3))}}));
  assign y5 = (3'd7);
  assign y6 = $unsigned({3{{4{b0}}}});
  assign y7 = (~^a2);
  assign y8 = (~{((!(~^b3))<<<(|{p12,p2,p16})),((~&{p7,p7})&{p1,p4})});
  assign y9 = (|(!((~&((b3?p5:b1)-(|p15)))<<(~(~&(p4>>>p12))))));
  assign y10 = {$unsigned(p5)};
  assign y11 = {$signed((b0+b1)),(~{3{b1}})};
  assign y12 = (5'd4);
  assign y13 = {{2{{b3,a3,b0}}},({a4,a2}!==$unsigned((a5>>>a0))),((b3?a1:b3)<<<(b1?a5:a1))};
  assign y14 = (~^({1{(+(~|{1{(b5-b5)}}))}}?($signed(b1)?(a3?a5:b5):(a0<<a2)):{4{{2{b4}}}}));
  assign y15 = (((b0!==b5)===(b5<<<b3))|{(p13!=p6),{(p7<<p7)}});
  assign y16 = (!{(b2===a2)});
  assign y17 = (~{4{(3'd6)}});
endmodule
