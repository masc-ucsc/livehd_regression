module expression_00013(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(5'd2 * (3'd4))}};
  localparam [4:0] p1 = (~&(+((5'd26)?(-5'sd15):(2'd0))));
  localparam [5:0] p2 = {(|({1{((-3'sd0)^~(3'd4))}}!=((4'sd1)^(4'sd6)))),(~|(~{2{{(~&(-2'sd1))}}}))};
  localparam signed [3:0] p3 = (!(&(((4'sd6)<<<(5'sd14))>={(3'd1),(2'd2),(5'd18)})));
  localparam signed [4:0] p4 = ((((4'd10)?(-5'sd9):(3'd5))?((4'd3)?(2'd1):(4'd15)):((-3'sd0)?(2'd1):(4'sd2)))?(-((4'd8)?(5'd16):(4'd11))):(|((5'sd13)?(5'sd4):(5'd6))));
  localparam signed [5:0] p5 = {1{(({4{(-5'sd14)}}?{3{(3'd7)}}:((-2'sd1)?(-2'sd0):(5'd16)))<=(((-5'sd13)-(5'd16))|{4{(-3'sd0)}}))}};
  localparam [3:0] p6 = ((({(2'd1)}^{2{(4'd9)}})&&{1{{(3'd5),(-5'sd5),(-3'sd3)}}})<=(({4{(3'd1)}}+((3'd3)<<<(2'd3)))&({(3'd1)}-((3'd1)|(4'd11)))));
  localparam [4:0] p7 = ((((3'sd3)-(3'd6))|{3{(4'd13)}})<<<(((3'd7)?(5'sd10):(3'd1))<<((-4'sd6)+(5'd9))));
  localparam [5:0] p8 = (((5'd10)!==(3'd3))%(-4'sd0));
  localparam signed [3:0] p9 = (((3'd5)?(3'sd3):(2'd1))|(&(2'sd0)));
  localparam signed [4:0] p10 = (4'd8);
  localparam signed [5:0] p11 = ((6'd2 * {3{(4'd5)}})===(((3'd0)!=(4'd14))&&((3'sd1)>=(-4'sd0))));
  localparam [3:0] p12 = (4'd14);
  localparam [4:0] p13 = {{(2'd3),(4'sd2),(-3'sd0)},((-3'sd2)?(5'd11):(4'd15))};
  localparam [5:0] p14 = (4'd4);
  localparam signed [3:0] p15 = (~(-((((-4'sd4)>>>(5'd23))===(-(-2'sd1)))>(((2'd2)!=(2'd0))&&((2'd3)&(3'd0))))));
  localparam signed [4:0] p16 = ((~&(-3'sd1))?((5'd27)*(5'sd13)):((2'sd0)?(3'd2):(5'sd15)));
  localparam signed [5:0] p17 = (-(2'd3));

  assign y0 = (({1{p4}}>>(b3?p16:a2))<<(-5'sd11));
  assign y1 = (((~a2)|{b4,b4,b2})^((b5!=b5)>>>(p10<=b0)));
  assign y2 = ({4{(-4'sd1)}}!==((((a3>>>b3)))>>>(-4'sd6)));
  assign y3 = ((~&((a2>>a1)>={4{a5}}))>>{2{(-b2)}});
  assign y4 = ($unsigned($unsigned((-3'sd0)))?((5'sd8)==$unsigned(p16)):$unsigned({a5,p0}));
  assign y5 = (b3|a2);
  assign y6 = ({((p8<a3)),{b3,b5,a3},((p9^b3))}>(((p7<<p12))|((b4)>>>{4{b1}})));
  assign y7 = {(b4&&b1),{p15}};
  assign y8 = $signed((-((|((!((b4===b4)>{(a1&&p17)}))))||(((b0<<b2)!==(|b0))<<{{p10,p17,p3}}))));
  assign y9 = (-(-(b4|a3)));
  assign y10 = (((p8&a0)|(2'd2))==((-3'sd3)||(2'sd0)));
  assign y11 = $unsigned({2{({4{p8}}?{3{a0}}:(-5'sd5))}});
  assign y12 = ((p2+b1)&&(b2>b4));
  assign y13 = ((((b0?b3:p14)&(b4?a3:p8))||((a5?b0:a0)^~(p9>p15)))+(-3'sd2));
  assign y14 = {2{{(b3===a0),{4{p10}},{2{p6}}}}};
  assign y15 = (p4==p3);
  assign y16 = (((~(-b4))<(&(p0!=p3)))<<<{3{{1{p1}}}});
  assign y17 = (3'd4);
endmodule
