module expression_00765(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~|((^((4'sd0)|(2'd3)))>>>(2'd0)))-(((5'sd3)?(3'd4):(4'sd2))!=((5'd6)^(3'd4))));
  localparam [4:0] p1 = (~|(5'sd11));
  localparam [5:0] p2 = ({3{(-4'sd7)}}<<(|(~&(4'd7))));
  localparam signed [3:0] p3 = (4'sd6);
  localparam signed [4:0] p4 = ((-2'sd0)?(!(5'sd0)):(4'd9));
  localparam signed [5:0] p5 = {4{(4'd9)}};
  localparam [3:0] p6 = (-3'sd3);
  localparam [4:0] p7 = ((6'd2 * ((4'd8)==(4'd1)))^{(5'sd3),(-2'sd1),(5'sd1)});
  localparam [5:0] p8 = {4{(3'sd2)}};
  localparam signed [3:0] p9 = (+((^((4'sd4)>(2'd3)))*(+(-4'sd4))));
  localparam signed [4:0] p10 = {1{{1{(~(({(2'd3),(2'd2)}^(~^(2'd0)))?{2{((-3'sd3)!==(2'sd1))}}:((3'd0)?(3'd7):(-5'sd12))))}}}};
  localparam signed [5:0] p11 = (5'd15);
  localparam [3:0] p12 = (~{1{(3'd2)}});
  localparam [4:0] p13 = (|(({(3'd4),(4'd14),(4'sd6)}?(~|(2'd3)):((3'd5)|(4'd15)))>>>{{(2'd1),(3'd7)},(!(3'd3)),(-3'sd0)}));
  localparam [5:0] p14 = (-2'sd0);
  localparam signed [3:0] p15 = (+(2'sd0));
  localparam signed [4:0] p16 = ({(3'd3),(2'd0),(-4'sd6)}?(~|(2'd2)):((-5'sd1)>>>(3'sd0)));
  localparam signed [5:0] p17 = (((5'd2 * (4'd5))>=((4'd11)^(3'd4)))?(((4'sd7)?(-4'sd5):(3'd6))|((5'd5)-(4'sd1))):(((-4'sd4)==(-4'sd5))?((-3'sd3)==(-4'sd3)):((5'd11)?(-2'sd0):(-4'sd2))));

  assign y0 = ((a1?b0:b2)?(3'sd0):(5'd11));
  assign y1 = {1{((^(!(a5===b1)))?((~b4)?(b1?b2:b4):(~b5)):((~|b1)?(a2?a0:a1):(b5?a1:p10)))}};
  assign y2 = ((-5'sd1)<={p1});
  assign y3 = {1{(-2'sd1)}};
  assign y4 = (a5!=b1);
  assign y5 = {(4'd4),$signed((^{(~^b3)}))};
  assign y6 = (2'sd0);
  assign y7 = (((-(-a3))<<(~|(a1+p9)))<<<(-{(a1?b4:a3),(b2?a1:b2),{a2,b0,a4}}));
  assign y8 = (p10+p17);
  assign y9 = (3'd6);
  assign y10 = ((2'd0)&&((a1!==b5)?(p6>>a0):(3'd2)));
  assign y11 = (^((2'sd1)|(b2&&a3)));
  assign y12 = ((a4!==b0)?(a4?b5:p11):(p8?p0:p7));
  assign y13 = {$unsigned((3'sd0))};
  assign y14 = {(b5?p12:p7),(b3)};
  assign y15 = {1{$signed({(p15),$unsigned(p0),(p15<<p0)})}};
  assign y16 = (~^$signed((-5'sd4)));
  assign y17 = (4'sd4);
endmodule
