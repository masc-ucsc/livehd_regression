module expression_00797(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-4'sd3)|((2'sd0)^~((4'd10)>(-2'sd0))));
  localparam [4:0] p1 = (~(!((((2'd2)?(4'sd4):(2'sd0))>((4'd12)!==(3'd2)))^(((5'd6)==(3'd4))-((3'd2)!=(3'd7))))));
  localparam [5:0] p2 = ((5'd2 * (4'd4))>(!(3'd5)));
  localparam signed [3:0] p3 = (((4'd11)^~(2'd0))&((-4'sd1)&(-4'sd7)));
  localparam signed [4:0] p4 = (~&({2{(|(-(3'd0)))}}||({2{(4'd6)}}<<((-4'sd0)^~(4'd8)))));
  localparam signed [5:0] p5 = (-(~|(3'sd2)));
  localparam [3:0] p6 = ((5'd5)?(-4'sd7):(5'd13));
  localparam [4:0] p7 = (((3'd5)|(-5'sd15))>={(-2'sd0),(5'd27)});
  localparam [5:0] p8 = (2'sd1);
  localparam signed [3:0] p9 = ((4'd0)<(5'd11));
  localparam signed [4:0] p10 = (2'd1);
  localparam signed [5:0] p11 = (((-5'sd12)===(3'sd2))/(3'd0));
  localparam [3:0] p12 = ((3'd5)%(5'sd5));
  localparam [4:0] p13 = (((3'd5)?(2'd1):(5'sd10))?{((2'd3)>(5'd18))}:(&((4'sd3)?(2'd2):(5'd3))));
  localparam [5:0] p14 = ({((4'd8)?(5'd21):(4'd0))}?{4{(2'd0)}}:{(!{4{(-3'sd2)}})});
  localparam signed [3:0] p15 = (-(~|((((3'sd0)>>(3'd5))>=((2'd2)^~(5'd22)))-(((3'd5)?(5'd26):(-4'sd6))===((5'd15)==(4'sd6))))));
  localparam signed [4:0] p16 = (((5'd2 * (4'd15))>((2'd0)>>>(4'd5)))|(((5'sd10)<<<(4'd4))^((2'd3)<<<(-4'sd3))));
  localparam signed [5:0] p17 = (-4'sd5);

  assign y0 = (4'sd5);
  assign y1 = {(((a4>>>a1)&{4{a4}})!=={(b1&a3),(a1>=b0)})};
  assign y2 = $signed((-5'sd0));
  assign y3 = $unsigned((5'd28));
  assign y4 = (3'd0);
  assign y5 = (!(~((~&(-(|b0)))^~{b2,b3,a2})));
  assign y6 = {{2{(~{p5,p6})}},{1{((p6<=b2)!=(p9&&p7))}},{2{{a4,b4}}}};
  assign y7 = {1{{2{(b1>=a2)}}}};
  assign y8 = {2{({3{(-2'sd0)}})}};
  assign y9 = (!{(|({4{b2}}?{p9,p17,b4}:(b0?p0:p7)))});
  assign y10 = $unsigned((((-5'sd4)*$signed((3'd6)))^~($unsigned((b1^~a0))==$signed((a4!=a3)))));
  assign y11 = (((a0?a3:b5)?(b3):(2'd1))?((6'd2 * b0)/b4):(((2'd1))<<(a4?b4:b5)));
  assign y12 = ((~&({(p6>=p12),(+p17)}<<((-p9)<<<(b3?a0:b2))))<((p16<p13)?(a0&b4):(p7<=p7)));
  assign y13 = ((5'sd12)<<<{(&p1),(a0<p10),(p0)});
  assign y14 = ((a2?a5:p8)>>>(b5>a2));
  assign y15 = $signed($unsigned(((~($signed((a0<b5))&(a3<b0)))<=$signed(((a2|b1)>(a1&&p15))))));
  assign y16 = (((3'd4)<<<(3'sd0))>(-3'sd2));
  assign y17 = ((a1>=a2)<=(b2===b1));
endmodule
