module expression_00995(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&(-((~^(5'd16))|(((3'd4)?(-5'sd0):(2'sd1))>>((-2'sd1)&&(4'd5))))));
  localparam [4:0] p1 = (((-2'sd0)?(5'd28):(-3'sd0))?((2'd3)?(3'sd2):(5'd19)):((4'sd1)?(3'd5):(3'd5)));
  localparam [5:0] p2 = (4'sd6);
  localparam signed [3:0] p3 = (5'd23);
  localparam signed [4:0] p4 = (~&(~^(2'sd0)));
  localparam signed [5:0] p5 = {4{(|(-2'sd1))}};
  localparam [3:0] p6 = (((2'd0)?(-((5'sd12)|(-5'sd14))):((2'd3)?(-2'sd1):(3'd6)))>>(5'sd10));
  localparam [4:0] p7 = ({2{(~&(-2'sd0))}}^{3{(3'sd1)}});
  localparam [5:0] p8 = ({((4'd9)-(4'sd0)),{(^(2'sd0))}}-(&{((5'd21)-(4'd15)),((-5'sd15)&(4'd9))}));
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = (~&{(~&(~|(-4'sd2))),{(5'd17),(2'd0),(2'sd0)},(|(&(2'sd1)))});
  localparam signed [5:0] p11 = ((!(~|{(2'sd1),(4'd9),(-4'sd4)}))>={((2'sd1)<=(-2'sd0)),{(5'd8),(-4'sd3),(2'sd1)}});
  localparam [3:0] p12 = {2{{((-4'sd2)&&(-5'sd15)),{3{(4'sd3)}},{1{(-5'sd6)}}}}};
  localparam [4:0] p13 = {(-(~(+(~^(^((-5'sd12)!==(3'd6)))))))};
  localparam [5:0] p14 = (~&(!(((5'sd12)?(-5'sd0):(5'd22))&(~|((5'd11)?(5'sd15):(2'd0))))));
  localparam signed [3:0] p15 = ((-3'sd3)?(~^(4'd4)):(3'd2));
  localparam signed [4:0] p16 = {3{(3'd7)}};
  localparam signed [5:0] p17 = ((5'd13)||(5'd16));

  assign y0 = (~&(a5^~b4));
  assign y1 = {{1{(a2==a4)}},(a5?p6:a0),(2'd1)};
  assign y2 = {($signed((&p1))?(p13^~a3):$signed((a0||a5))),({$unsigned(b4),(-a0)}<=$unsigned((p6>>b0)))};
  assign y3 = (((a0?p7:p11)>>>(p3%a5))?(p16?p4:p6):(p15?p1:p6));
  assign y4 = {(b2<=p3),{p12,p12},{b0,p16,p4}};
  assign y5 = (&(~&$unsigned((!(3'd6)))));
  assign y6 = ({3{p10}}?(a5!==b3):(a5?b5:p15));
  assign y7 = ((b2?p9:b0)?(a3?a5:b4):(b2&a0));
  assign y8 = {3{(((p5?p14:a2)))}};
  assign y9 = (~^(!((a4?b2:b0)?$signed((!(|a5))):(+$signed((a0))))));
  assign y10 = {p8,p12,a1};
  assign y11 = (&({{p13},(-b3)}?({b2}<(p1|a5)):(&{p12,a3,p6})));
  assign y12 = ({(b0)}?(b1==a1):(p5|b1));
  assign y13 = $signed((4'd2 * (^(4'd9))));
  assign y14 = (+{4{{3{p0}}}});
  assign y15 = ({({p16}<(5'd29))});
  assign y16 = ((3'sd2)>>((6'd2 * b2)?(a0?a2:a5):(6'd2 * b1)));
  assign y17 = {(~|{(&(~&(&a5))),(|(-{p2}))})};
endmodule
