module expression_00183(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(3'd6));
  localparam [4:0] p1 = (&(5'd19));
  localparam [5:0] p2 = {{{(2'd3)}}};
  localparam signed [3:0] p3 = (^{3{(~&(5'd2 * (5'd18)))}});
  localparam signed [4:0] p4 = (2'd0);
  localparam signed [5:0] p5 = ({4{(-5'sd14)}}-{4{{1{(4'd7)}}}});
  localparam [3:0] p6 = ({(-2'sd0),(4'd13)}?(|(5'd2)):(~|(5'sd2)));
  localparam [4:0] p7 = {{(2'd1),(2'd2),(3'd7)},((5'd17)>=(4'sd7)),((-2'sd0)==(3'd0))};
  localparam [5:0] p8 = (((4'd8)<=(3'd4))-((4'sd7)>>>(2'd3)));
  localparam signed [3:0] p9 = ((-4'sd6)?(2'd0):(2'd2));
  localparam signed [4:0] p10 = ((4'd4)|(5'd15));
  localparam signed [5:0] p11 = (((2'd2)&(3'd1))>>>((3'sd2)|(-3'sd2)));
  localparam [3:0] p12 = ({{(5'd13),(4'sd0)},((5'sd15)===(4'd9))}<{3{((2'd3)!=(-3'sd3))}});
  localparam [4:0] p13 = (4'd2 * (!(~^(3'd5))));
  localparam [5:0] p14 = ((~^((2'd3)?(-4'sd3):(-5'sd8)))?(|((!(2'd2))&&((5'sd12)?(3'd0):(-2'sd0)))):(+((-(3'd2))^~((2'd3)?(2'd3):(4'sd7)))));
  localparam signed [3:0] p15 = (+{3{(4'd1)}});
  localparam signed [4:0] p16 = (-4'sd3);
  localparam signed [5:0] p17 = (-2'sd0);

  assign y0 = (((a1?p2:b1)/a0)>=(~(((a0%a3)>(b1||p11))-(a4?b3:p13))));
  assign y1 = {4{{1{(&(~|$unsigned(p16)))}}}};
  assign y2 = (((b5+p2)?(a4?p12:p10):(^(b0===b3)))>>>(((!p1)>>>(5'sd1))|((~^p10)||(p14?a0:p7))));
  assign y3 = (({b5,a5}?(b5?a5:b2):{a1,a1})?$unsigned({{a0},{a3,a1}}):{{b2,a3},{p0},{a2,p3,a0}});
  assign y4 = ({1{(^(((b2+b2)<<{1{a5}})|((b4?b2:b2)||(a2!==a0))))}}===(5'd2 * (a0<<<b2)));
  assign y5 = ($signed({3{a1}})<<<(&(b0|p0)));
  assign y6 = ((a2?a1:a3)!==(a5?b3:b3));
  assign y7 = {(b0===b3),(b3>>a0),{b5}};
  assign y8 = {3{p14}};
  assign y9 = {2{(((a4<<p16)<<<(p0)))}};
  assign y10 = (!{4{(~a2)}});
  assign y11 = (((b1|a3)!=(b2===b1))||{1{(a1===a1)}});
  assign y12 = (p7^b0);
  assign y13 = {$unsigned(b0),{1{p13}},(^b0)};
  assign y14 = {b3,a3};
  assign y15 = {1{(~&((((p0>>p11)|(~|$unsigned(p3))))>$signed({1{(6'd2 * $unsigned((b3===a2)))}})))}};
  assign y16 = {1{(~|(p13|b4))}};
  assign y17 = {$unsigned(($unsigned((!{{4{a0}}}))>={4{(p12)}}))};
endmodule
