module expression_00502(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-5'sd0);
  localparam [4:0] p1 = (~{(5'd15),(-5'sd12)});
  localparam [5:0] p2 = (-(~^((+(~|(~^(3'd6))))!=(&(~^((2'd3)?(2'd2):(-4'sd7)))))));
  localparam signed [3:0] p3 = ((3'd2)>>>({2{(2'sd1)}}>>(5'd22)));
  localparam signed [4:0] p4 = {1{(5'sd9)}};
  localparam signed [5:0] p5 = (+(({1{{1{(4'sd7)}}}}>=(~|{3{(5'd20)}}))||({1{{4{(-3'sd1)}}}}<<<(-{3{(-3'sd3)}}))));
  localparam [3:0] p6 = ((~^(-{(-((4'sd6)^~(-3'sd1)))}))<<(-{((5'd22)||(4'sd7)),(^(5'd6)),((3'd7)?(4'd2):(4'sd1))}));
  localparam [4:0] p7 = (^(5'd11));
  localparam [5:0] p8 = (&{{(4'd3),(-2'sd0)}});
  localparam signed [3:0] p9 = (+(~&(3'd7)));
  localparam signed [4:0] p10 = ((-5'sd0)>>>(5'd26));
  localparam signed [5:0] p11 = ((~&(|((!(3'sd0))?((3'sd0)?(2'd1):(3'sd1)):((3'sd1)<=(4'sd7)))))>(-5'sd4));
  localparam [3:0] p12 = ((4'sd3)===(2'd3));
  localparam [4:0] p13 = {4{(~^{{(-2'sd1),(5'd23),(-2'sd1)}})}};
  localparam [5:0] p14 = ((+(5'd25))===((4'sd1)==(3'd0)));
  localparam signed [3:0] p15 = (^(-{{{(~(-2'sd1)),(-(3'sd0)),(|(2'd0))}},{(~&(~|(~^{(2'sd1),(4'sd4),(4'sd2)})))}}));
  localparam signed [4:0] p16 = (((5'd14)?(-4'sd5):(3'd5))?(!(3'd2)):((2'd2)-(-4'sd1)));
  localparam signed [5:0] p17 = (((4'd6)^~(-4'sd3))>>>{(3'd7),(3'd7),(2'sd1)});

  assign y0 = (3'd3);
  assign y1 = {4{(p7&p8)}};
  assign y2 = {3{{b4}}};
  assign y3 = ((p2?a0:a1)!=(b4+b0));
  assign y4 = {((~$unsigned((+($signed(($unsigned(b1)<<<{b3,p11})))))))};
  assign y5 = (-(~{(-(a3?p10:p0)),{(+(p5!=p7))},((|p7)&(|p10))}));
  assign y6 = {4{($signed(a0)?(p6<<p17):{2{p11}})}};
  assign y7 = ((~(-5'sd13))?{{{a3},(p6>>p1)}}:((a2?b5:a3)<<<(5'd28)));
  assign y8 = {3{(!((+(b1|a5))<=(p8>>>b1)))}};
  assign y9 = (2'sd0);
  assign y10 = {3{$signed(({2{(5'd2 * b0)}}))}};
  assign y11 = {4{{3{p10}}}};
  assign y12 = ((a1?b4:b0)>(b2?a2:b5));
  assign y13 = (~^(a4||p9));
  assign y14 = ((({b1}^(~a5))^((a3==a3)^{2{a1}}))!=={1{{(~(b4&a1)),(4'd2 * {b2,b2})}}});
  assign y15 = (^{((b4?a1:p15)>=(p16)),(p12?p7:b0),($unsigned(a0)===(^a3))});
  assign y16 = {4{((a5?p6:p17)?{2{p2}}:{3{p11}})}};
  assign y17 = {(p14),(5'd2 * a0),(a0<=p0)};
endmodule
