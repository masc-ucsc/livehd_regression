module expression_00355(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{((~(-5'sd11))>(~(-5'sd12)))}};
  localparam [4:0] p1 = ({(3'd1),(3'd4),(-3'sd2)}<(3'd4));
  localparam [5:0] p2 = (|((+(~^{3{(-4'sd0)}}))>=(!{3{(3'd4)}})));
  localparam signed [3:0] p3 = ({(-2'sd1),(5'd31)}>>{(3'sd2),(-4'sd6)});
  localparam signed [4:0] p4 = (((4'd8)>=(-3'sd2))>((-3'sd0)!==(3'sd2)));
  localparam signed [5:0] p5 = (-3'sd3);
  localparam [3:0] p6 = ((((5'd26)?(3'd1):(3'sd2))?((3'd0)?(2'd2):(2'd3)):((-3'sd1)?(-2'sd0):(3'd7)))?(((-4'sd6)?(5'd24):(-5'sd8))?((3'd6)?(4'sd6):(-4'sd2)):((4'd7)?(5'd9):(-3'sd1))):(((5'd16)?(4'd2):(-5'sd13))?((-5'sd9)?(-4'sd6):(3'd7)):((4'sd0)?(2'sd1):(-2'sd1))));
  localparam [4:0] p7 = (-3'sd3);
  localparam [5:0] p8 = (((5'd23)?(-4'sd1):(-5'sd13))/(-2'sd0));
  localparam signed [3:0] p9 = (&(3'sd1));
  localparam signed [4:0] p10 = ((((5'd8)===(4'd11))?((4'sd7)?(5'd20):(5'd3)):{(5'sd5),(5'sd9)})>>(((2'd3)&(3'd0))===((-5'sd8)?(-4'sd4):(4'd15))));
  localparam signed [5:0] p11 = {3{{3{(-5'sd4)}}}};
  localparam [3:0] p12 = (((5'sd5)?(4'd10):(-4'sd4))?{(5'd15),(3'd3)}:((5'sd14)?(4'd10):(-4'sd7)));
  localparam [4:0] p13 = (^(2'd0));
  localparam [5:0] p14 = (~&(^(3'd4)));
  localparam signed [3:0] p15 = {1{(~{1{(~&(3'd6))}})}};
  localparam signed [4:0] p16 = (^(!({((2'sd0)<<(2'sd0)),{(5'sd0),(4'd5)}}+(~^((-(3'sd2))!=((4'd3)+(-4'sd0)))))));
  localparam signed [5:0] p17 = (5'd17);

  assign y0 = (((b4&b5)>{b5})===(!{4{a1}}));
  assign y1 = ($signed((~^$unsigned($unsigned((((~^b5)&&$signed(a3)))))))!==((^((a5||b4)&&(b3<<<b5)))));
  assign y2 = (({b5,a4}?(b2<<<a3):(b3?b1:b0))?{((p0?b3:b1)?(b0?p17:a0):{a1,a0,p14})}:({(p0?a0:b0)}>(a5===b3)));
  assign y3 = (a1||b5);
  assign y4 = ((5'sd13)?(&({2{p13}})):(5'd2 * (p12?b0:p7)));
  assign y5 = ((|((a3?b5:b0)/a4))>>(|(&((-(a3+a2))?(!(+p0)):(b3?b0:a1)))));
  assign y6 = ({({p14,p14}&&(p11>p6))}<=(((p5>=p13)<<<(p1^p16))<={(p7<=p6)}));
  assign y7 = ((b0>a3)?(b1!==a1):(-p16));
  assign y8 = {2{(a1+a4)}};
  assign y9 = (~($signed((!(|({2{b5}}<{2{a4}}))))>(((a4^b3)^~(p11^b4))&&($unsigned(b0)&(~a1)))));
  assign y10 = {2{((p2>=p7)+{p8,a2})}};
  assign y11 = ($signed({$unsigned((b2^b3)),$signed((p12<=p5))}));
  assign y12 = (~^$unsigned(({4{p11}}=={1{{2{p1}}}})));
  assign y13 = (|((4'd6)^(^((b2<b2)/a2))));
  assign y14 = (5'sd6);
  assign y15 = {4{(~|{1{p14}})}};
  assign y16 = (!(~&((^(p13/p15))||(~|(!(~^b5))))));
  assign y17 = ((-{1{((6'd2 * (b0>>b2))>>>{3{a4}})}})^~{4{(a1<=b3)}});
endmodule
