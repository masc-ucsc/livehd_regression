module expression_00265(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(~((-3'sd3)?(2'd1):((2'd0)+(5'd15)))));
  localparam [4:0] p1 = (-2'sd1);
  localparam [5:0] p2 = ((4'd9)?(2'd1):(-3'sd3));
  localparam signed [3:0] p3 = ((((3'd0)?(3'd0):(3'sd3))>>((5'd15)^~(-5'sd8)))?(((4'd5)?(3'd0):(5'd9))>((5'd8)?(2'd3):(-5'sd14))):{{2{(2'sd0)}}});
  localparam signed [4:0] p4 = {{(-4'sd6)},((5'd8)|(2'd1)),{(4'sd2)}};
  localparam signed [5:0] p5 = (^((|(4'd4))<=((4'd14)==(4'd3))));
  localparam [3:0] p6 = (|(^(5'd2 * (-(~&(2'd0))))));
  localparam [4:0] p7 = {(-4'sd0)};
  localparam [5:0] p8 = ({1{{((4'sd4)&(2'd1)),((3'd1)&(2'd3)),{(3'd2),(5'd30)}}}}!==(|({4{(2'sd0)}}&&(+(4'd0)))));
  localparam signed [3:0] p9 = ({1{(6'd2 * ((4'd3)<(4'd11)))}}>(^{(5'd2 * (2'd0))}));
  localparam signed [4:0] p10 = {(~&{(3'd0)}),(-{(4'd4)})};
  localparam signed [5:0] p11 = ((~&(~{4{(2'd3)}}))>={2{((2'sd1)<<<(2'sd0))}});
  localparam [3:0] p12 = (5'd8);
  localparam [4:0] p13 = (~&((((5'sd9)<(4'd12))==={1{(4'd3)}})>>>{4{(3'd6)}}));
  localparam [5:0] p14 = ((3'd5)>>(4'd15));
  localparam signed [3:0] p15 = ((-4'sd4)<=(-5'sd9));
  localparam signed [4:0] p16 = {{(-5'sd13),(-4'sd0)},{(-2'sd0),(-3'sd0),(-2'sd1)},((3'd1)<<<(4'd6))};
  localparam signed [5:0] p17 = ({3{(4'd5)}}==={4{(4'sd6)}});

  assign y0 = ((&{{a1,b3,b1}})>>>({p6,a2}-(!{b3,b4})));
  assign y1 = (($unsigned(p4)&{3{b1}})>>(3'd2));
  assign y2 = (a1?b3:a1);
  assign y3 = {3{(4'sd0)}};
  assign y4 = ({p12,p14}-(~&p13));
  assign y5 = (((p4?p8:a3)^~(3'sd3))?((~|(b5!==a0))|(-3'sd3)):({3{b5}}!==(&(4'd13))));
  assign y6 = (^$signed($signed($signed(p2))));
  assign y7 = (((|$signed(p16))/p16)==((6'd2 * (+$unsigned(p15)))<(!((p6||p4)&&(p16<<p17)))));
  assign y8 = (~|(-(~&{3{p13}})));
  assign y9 = (~|((p14>>b1)/a3));
  assign y10 = ({3{(a2<<a5)}}!==((3'd3)));
  assign y11 = {{(p14>p9),(5'sd10)},((3'd5)<<{p15,a4,p11}),(2'd2)};
  assign y12 = (3'd2);
  assign y13 = {(~^({(b2<<<a3),(a2<p16),(p4<<a5)}&(!(~^(~(&(~&b2)))))))};
  assign y14 = $unsigned(((((-(+(b4|a4)))+(~&{1{(b4<<b0)}})))&&(((b3|b4)||(~&a4))<=({1{p10}}>>>{2{a0}}))));
  assign y15 = (~|(~^(-(&(-4'sd4)))));
  assign y16 = ((b0?b1:a0));
  assign y17 = ({1{{1{{2{$signed({1{{4{p9}}}})}}}}}});
endmodule
