module expression_00837(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(|(((5'sd8)||(3'sd1))^(~{(4'sd0)}))));
  localparam [4:0] p1 = {4{((2'sd0)?(5'd7):(3'd0))}};
  localparam [5:0] p2 = (((!(2'sd0))<=((-3'sd1)<<<(-4'sd3)))|{((~&(5'sd8))|((5'd14)<(-4'sd7)))});
  localparam signed [3:0] p3 = ((3'd3)-(2'd2));
  localparam signed [4:0] p4 = {(-4'sd2),(3'd5)};
  localparam signed [5:0] p5 = (({3{(4'sd5)}}?(-(-5'sd15)):((2'sd0)?(2'sd1):(3'd5)))&((|((2'd2)<(5'd24)))>((-5'sd3)>>(4'sd6))));
  localparam [3:0] p6 = (~&{2{(~|(+(2'd0)))}});
  localparam [4:0] p7 = ((-3'sd1)?(!((-3'sd2)?(3'd4):(-3'sd3))):(5'd18));
  localparam [5:0] p8 = {(((4'd14)?(4'sd6):(4'd3))<(-{((3'sd3)&&(-5'sd13))})),(&((^((5'sd5)?(-2'sd0):(3'd2)))>>{(3'd0),(3'd5)}))};
  localparam signed [3:0] p9 = {2{(4'sd7)}};
  localparam signed [4:0] p10 = {1{(~&(({4{(4'sd3)}}-((3'sd1)<(-3'sd2)))&&({4{(5'd29)}}||(4'd2 * (5'd18)))))}};
  localparam signed [5:0] p11 = (((-2'sd0)^~(2'd1))||{(-2'sd0),(5'd27),(5'd5)});
  localparam [3:0] p12 = (((5'd5)?(-5'sd6):(3'sd2))?((5'sd1)%(4'd3)):((2'd1)?(3'd5):(-3'sd3)));
  localparam [4:0] p13 = ((-(-((5'sd5)?(5'd4):(3'd1))))>=(&{2{(5'sd10)}}));
  localparam [5:0] p14 = {{(4'd5),(3'd6),(3'd3)},{(-5'sd3)}};
  localparam signed [3:0] p15 = (-(5'd5));
  localparam signed [4:0] p16 = ((5'd9)?(3'd6):(-3'sd3));
  localparam signed [5:0] p17 = {2{(4'd2)}};

  assign y0 = (((b1?b0:b5)|{a1,a4,b2})!==({b1,b5}?(a5|a0):{2{b0}}));
  assign y1 = {4{(&(p3^~b3))}};
  assign y2 = (~^{3{{1{(+b5)}}}});
  assign y3 = (p3?p3:p8);
  assign y4 = (5'd7);
  assign y5 = (^{1{({{(b3>p6),(a1^~a3)}}<<<({3{p14}}^~(b3===a2)))}});
  assign y6 = (6'd2 * (4'd12));
  assign y7 = (p3&&b0);
  assign y8 = ((+(|p14))==(~(~p15)));
  assign y9 = (+((2'sd1)?((a4?a3:b4)?(a1?b0:b5):(a4?a5:p14)):(-4'sd3)));
  assign y10 = ((+(p8?a0:a4))||{b4,b1});
  assign y11 = (3'd1);
  assign y12 = $signed(({1{$signed((5'd9))}}));
  assign y13 = $signed(($unsigned((p7>>>p11))+(^$unsigned(p3))));
  assign y14 = {1{{2{({3{p13}}?(p12?p8:p1):(p8<<p11))}}}};
  assign y15 = {{p1,p2},(^p7)};
  assign y16 = ({(a0?b1:p7),(b2?b5:p3)}?$unsigned((p7?p3:p12)):{p5,p15,p13});
  assign y17 = ((-(~^p10))*(+(p15-p1)));
endmodule
