module expression_00537(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((|(~^(~|(^(5'd7)))))^(~^(((4'd14)!==(-2'sd0))/(-2'sd1))));
  localparam [4:0] p1 = ((((3'd2)>>>(3'd2))/(5'd26))^(((4'd7)*(5'sd10))|(~&((4'd9)|(2'd0)))));
  localparam [5:0] p2 = (5'd2);
  localparam signed [3:0] p3 = (((-2'sd0)&&(2'd2))-((-4'sd4)&(-5'sd14)));
  localparam signed [4:0] p4 = ((&{(-3'sd0),(-4'sd7)})+((4'd2)?(2'sd1):(-5'sd0)));
  localparam signed [5:0] p5 = ({(!((2'd1)?(5'd8):(2'sd1))),(((3'd6)?(4'sd0):(-2'sd1))>={(5'd22)})}-(((4'd7)?(-5'sd14):(4'd6))?{((2'sd0)?(3'd1):(2'd3))}:(~|{(-4'sd3),(2'd0),(-2'sd1)})));
  localparam [3:0] p6 = {{(2'd2),(3'd6)},((2'sd0)-(2'sd1)),(4'd2 * (4'd6))};
  localparam [4:0] p7 = (((4'd4)<(3'sd1))|(-3'sd1));
  localparam [5:0] p8 = (({1{((3'sd1)<<(-5'sd2))}}-{((5'd30)==(2'd2))})<<(((-3'sd0)&&(4'd11))^~((-2'sd1)-(-2'sd0))));
  localparam signed [3:0] p9 = ((((3'd2)%(2'd3))+((2'd2)*(2'sd0)))?(((5'sd4)==(-5'sd12))>>>((5'd19)<=(4'd15))):(~|(&((5'd20)?(4'sd2):(-5'sd15)))));
  localparam signed [4:0] p10 = ((-3'sd1)&(2'sd0));
  localparam signed [5:0] p11 = {{4{(-3'sd1)}},{{2{{(-3'sd3),(-5'sd11)}}}}};
  localparam [3:0] p12 = (({4{(4'd6)}}&(!(-3'sd1)))!=(((2'd1)>>>(4'd1))<<<((-3'sd3)>=(-4'sd6))));
  localparam [4:0] p13 = (((5'sd0)!==((-4'sd5)==(2'd1)))?(2'd3):((3'sd2)?((4'd9)||(5'sd1)):((5'd2)?(4'd13):(2'sd0))));
  localparam [5:0] p14 = (((5'd21)<=(-3'sd2))>>>((5'sd9)>>>(3'd1)));
  localparam signed [3:0] p15 = {(-3'sd3),(2'sd1),(5'd17)};
  localparam signed [4:0] p16 = (((((3'd7)==(4'sd6))&{(5'd29),(-2'sd0)})=={(~&(-5'sd12)),((-5'sd13)&(-3'sd1))})!=={(&(&(4'd7))),((4'd4)<(5'd17)),((-5'sd5)===(5'd11))});
  localparam signed [5:0] p17 = {{((-5'sd8)<(4'd7)),{4{(4'd0)}},((4'd8)<=(4'd12))},(((4'd10)?(3'sd3):(2'sd1))?{(3'd2)}:((4'd5)?(-5'sd13):(2'd2)))};

  assign y0 = ($signed(p1));
  assign y1 = {3{{4{{1{p0}}}}}};
  assign y2 = ((~^((+b5)>>(a2!=a1)))^((~|a5)<<<(-p9)));
  assign y3 = {(~&(~^{(!(4'd2 * $unsigned(b0))),((~|a4)|(a0?a2:b1)),((b0!==b4)?(a4-a2):{a1,a1,b2})}))};
  assign y4 = ((6'd2 * b1)===(-2'sd0));
  assign y5 = (-(|((&$signed(p6))&(~^(5'sd10)))));
  assign y6 = (({(~|p15)}>={b1,p17})&&{$unsigned({p9,p10,p5}),(~^(a3||p3))});
  assign y7 = (a4|a0);
  assign y8 = {((a3?a1:b0)&&(b5-a0)),((p8^b3)?{p10}:(p3|b0))};
  assign y9 = (!$unsigned(({3{a0}}?(b2<<b5):{1{{3{a1}}}})));
  assign y10 = {2{(6'd2 * (a0?p12:p2))}};
  assign y11 = (((-4'sd3)&&(b4?p15:b3))?{(b4<p16),(p15?p11:b0),(&b1)}:(-4'sd6));
  assign y12 = (((2'd2)>=$signed((p2^p14)))!=(((p1^~p0)!=(p16))));
  assign y13 = (5'sd7);
  assign y14 = {({(p11&&b1)}),((p6)>(~^p2)),((^a5)>>>(p11==a4))};
  assign y15 = (^((!((~|b3)))!==(b5?b4:a0)));
  assign y16 = (((b3<=p8)&&(!(a2>a3)))+(!((a4<a1)+(a3&&p12))));
  assign y17 = $signed($unsigned((((p8?p8:b3))?(5'd0):(b4^~p6))));
endmodule
