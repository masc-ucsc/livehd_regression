module expression_00918(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|((~(((5'd5)&&(-2'sd1))||(!(2'sd0))))>>((-(5'sd11))<((2'd2)*(-4'sd4)))));
  localparam [4:0] p1 = {4{(&(^((-2'sd0)?(4'd1):(4'sd1))))}};
  localparam [5:0] p2 = ((((5'd27)>(-5'sd4))!==((-5'sd8)&(-4'sd2)))>>(((2'sd1)===(3'sd2))>>((3'd6)<=(3'd5))));
  localparam signed [3:0] p3 = ((((5'sd5)>(3'd1))|((3'sd1)&&(3'd0)))>({4{(5'd24)}}<<((3'd3)?(5'd0):(3'd5))));
  localparam signed [4:0] p4 = ({4{(5'd2 * (2'd0))}}+{3{(&(5'd13))}});
  localparam signed [5:0] p5 = (((3'sd1)!=(4'd8))<<<{4{(2'd3)}});
  localparam [3:0] p6 = ((-4'sd7)?(3'd7):(3'd5));
  localparam [4:0] p7 = ((+((4'd1)?(-2'sd1):(3'sd0)))?(!((3'd2)?(5'd26):(2'd1))):(|((3'sd2)?(3'd5):(-2'sd0))));
  localparam [5:0] p8 = (-3'sd2);
  localparam signed [3:0] p9 = {3{(4'd5)}};
  localparam signed [4:0] p10 = ((((4'd14)?(4'd7):(2'd0))?(2'd0):((3'sd3)<<<(4'sd5)))-(-2'sd0));
  localparam signed [5:0] p11 = (2'd0);
  localparam [3:0] p12 = (~&(!((((3'd4)==(-5'sd14))|(+(~&(-2'sd0))))!=((&(|(-4'sd3)))<=(~((-4'sd1)+(-4'sd3)))))));
  localparam [4:0] p13 = ((3'd5)!=(2'sd0));
  localparam [5:0] p14 = (~{(4'sd3),{3{(4'd3)}}});
  localparam signed [3:0] p15 = (!((~|((-2'sd0)>>>(-2'sd0)))<{((3'sd0)?(4'd8):(2'sd0)),{(5'd21),(3'sd2),(-3'sd3)}}));
  localparam signed [4:0] p16 = (-(3'sd2));
  localparam signed [5:0] p17 = {4{((2'd1)?(-2'sd0):(4'sd4))}};

  assign y0 = $unsigned((b0||p15));
  assign y1 = ((p4?p16:p3)?{4{p3}}:{3{p5}});
  assign y2 = ((^b4)-(5'd2 * b0));
  assign y3 = (3'sd2);
  assign y4 = {3{(a2==a5)}};
  assign y5 = {(5'd12)};
  assign y6 = {1{{2{(b0?a0:a5)}}}};
  assign y7 = ((3'sd2)>=(5'd6));
  assign y8 = (-5'sd11);
  assign y9 = (((p8<p16)||(p8^~p10))==((p4?p1:p13)?(p17<=p13):(p9<<<p10)));
  assign y10 = $unsigned({(!((|p17)<<(~p8))),$unsigned((&(3'd2))),{(p3?a3:a5),{b4,b3},{p11,a0}}});
  assign y11 = (5'd22);
  assign y12 = (6'd2 * p8);
  assign y13 = {$unsigned($unsigned((((p5?a1:a2))?{{b0}}:{{a5,a4}})))};
  assign y14 = (2'sd1);
  assign y15 = ((b4?p15:p2)-(a2?p7:p9));
  assign y16 = ((({b5}^(b1-b1))^((b1<<p0)|(b0?a5:a0))));
  assign y17 = {4{((p16&&p10)>>>(a4===b0))}};
endmodule
