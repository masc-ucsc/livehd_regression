module expression_00452(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-4'sd3)===(3'd1));
  localparam [4:0] p1 = {((5'd2 * ((3'd5)>>>(3'd1)))!=({(-3'sd2),(5'd20),(-4'sd4)}?{(2'd3),(5'd23),(4'd15)}:((3'd4)<<<(4'd10))))};
  localparam [5:0] p2 = ((3'd4)<<<(~&{2{(-5'sd10)}}));
  localparam signed [3:0] p3 = (~&(~&(~&{2{{2{((2'd1)===(4'd15))}}}})));
  localparam signed [4:0] p4 = (((5'sd8)|(-2'sd1))%(4'd4));
  localparam signed [5:0] p5 = ((&(+(((-3'sd1)==(-2'sd0))?((5'd20)&&(4'd6)):((3'd4)?(-3'sd2):(5'd11)))))<=(((5'd13)-(5'sd9))?(|((3'd3)===(4'd8))):(!((5'sd2)>>>(4'd7)))));
  localparam [3:0] p6 = (+((5'd24)<(3'd7)));
  localparam [4:0] p7 = {2{(((3'd2)>>>(5'd2))!=((-5'sd5)!=(2'd3)))}};
  localparam [5:0] p8 = ((((-5'sd10)?(2'd0):(4'sd7))>>((2'd3)?(2'd0):(4'd14)))>>>(((4'd13)?(2'd0):(2'd3))<<(~&(4'd4))));
  localparam signed [3:0] p9 = {{4{(2'sd1)}},((4'sd6)?(3'd4):(-5'sd10)),{4{(5'sd4)}}};
  localparam signed [4:0] p10 = (^{(3'd4),(3'sd1)});
  localparam signed [5:0] p11 = (+((((-2'sd1)?(-3'sd0):(5'sd7))?((3'd5)|(-3'sd1)):((-2'sd0)<<<(5'd22)))^(((4'd2)?(5'd19):(2'd0))<{(5'sd5),(-4'sd7)})));
  localparam [3:0] p12 = (-(+(|({((2'd2)^~(2'd2)),{(-5'sd4)}}?(&(~|{(3'd0),(4'd11),(-3'sd2)})):((5'sd14)?(5'sd6):(-4'sd7))))));
  localparam [4:0] p13 = (({(-3'sd1),(5'sd2)}<<<(+(3'sd3)))&&(((2'd0)^~(-3'sd3))>>>((5'd20)^~(4'd4))));
  localparam [5:0] p14 = ({4{((4'd5)&(2'sd0))}}^{3{((-3'sd1)-(2'sd1))}});
  localparam signed [3:0] p15 = (((-4'sd2)?(2'd3):(5'd25))<<((4'd2)>=(-4'sd6)));
  localparam signed [4:0] p16 = (^(5'sd6));
  localparam signed [5:0] p17 = {(~|(5'd18)),(5'd21),(-(4'd0))};

  assign y0 = (($unsigned((^((p8?p13:p4))))));
  assign y1 = (((~(3'd6))<(-4'sd0))<<<($signed($signed(b0))^~$signed((~&b2))));
  assign y2 = (!(6'd2 * (-(~|a0))));
  assign y3 = (((b4!==a1)!=(+(p12<=p5)))||(~|($unsigned(p1)<(a4<p1))));
  assign y4 = ({2{(p15?p12:p15)}}^((a2===b4)+(p6||p4)));
  assign y5 = {1{((a1?a2:p10)?(2'd3):(~|(+{3{p14}})))}};
  assign y6 = {1{(&({1{(3'd0)}}&(|(((3'd3)^~{1{b5}})>=((p2<=a4)^(b2>b1))))))}};
  assign y7 = (((p14!=b5)?(a2&&p7):(b0>>p2))?((p2)?(p12?p2:p1):(p15&&b5)):($signed(p14)-(p14?a4:b2)));
  assign y8 = $signed((|{p0,p1,p5}));
  assign y9 = (((a0!==a1))^~($signed({p3})));
  assign y10 = {3{((p4?p14:p14)>(3'd4))}};
  assign y11 = (($unsigned(p11)?(-2'sd0):(p0<=p0))>>>$signed((($unsigned(p4))>(p17?p11:p6))));
  assign y12 = {4{b1}};
  assign y13 = (({p0,b0}<<{p9,p17,p9})-{(p3==b3)});
  assign y14 = ((($unsigned((a2%a2))/p8)>(-(&(~|(|$signed((~(b1>>>b3)))))))));
  assign y15 = ((($unsigned(p17)>(p8/a3))^~((p12?p1:p0)<=(4'd2 * p2)))^~(2'sd1));
  assign y16 = {2{a4}};
  assign y17 = ((p13<<p8)?(p14-p11):(p14>p17));
endmodule
