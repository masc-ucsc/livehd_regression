module expression_00204(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'sd2)>>(-4'sd5))>((2'd0)<<<(3'd6)))?(~^(|(~((-4'sd3)^(3'd0))))):(~|{1{((5'sd5)==(3'd2))}}));
  localparam [4:0] p1 = (|(3'd6));
  localparam [5:0] p2 = {{(^(4'sd7)),(~(5'd29))},{(4'd12),(3'd6),(2'd2)},{{{(4'd6),(4'd9),(2'd3)}}}};
  localparam signed [3:0] p3 = ((~&((5'sd10)>>(3'sd1)))*(4'd2 * (2'd1)));
  localparam signed [4:0] p4 = ((((4'd8)>>>(5'sd10))===((2'sd0)<<(2'd0)))^~{2{((-2'sd1)>=(4'd2))}});
  localparam signed [5:0] p5 = (((2'd1)>=(-5'sd0))?((+(2'd0))^(|(4'sd2))):(-2'sd0));
  localparam [3:0] p6 = (|(~^(2'd0)));
  localparam [4:0] p7 = (~&(((-2'sd0)==(-4'sd4))%(2'd2)));
  localparam [5:0] p8 = (4'd2 * (2'd1));
  localparam signed [3:0] p9 = ({(5'sd15),(2'd3)}|(^(5'd24)));
  localparam signed [4:0] p10 = {(~^{(+(-{(3'd6),(-2'sd0)})),{(&(2'd3)),(^(3'd5))}})};
  localparam signed [5:0] p11 = (-4'sd0);
  localparam [3:0] p12 = {{((3'd3)<=(-3'sd2)),((5'd9)==(5'sd15))},({(3'd1)}==={(5'd12),(3'd0),(3'd6)})};
  localparam [4:0] p13 = (5'd8);
  localparam [5:0] p14 = ((4'd2)!==(((2'd2)?(2'sd0):(-5'sd7))?((-3'sd2)<<(2'd2)):((-4'sd6)?(2'd1):(3'sd3))));
  localparam signed [3:0] p15 = (((-3'sd1)-(5'd4))/(3'd6));
  localparam signed [4:0] p16 = (((3'sd0)!=(5'd30))?((-5'sd3)>>(-3'sd0)):((-5'sd0)?(-4'sd1):(-2'sd0)));
  localparam signed [5:0] p17 = ((((-2'sd1)<<<(5'd14))>=(!(2'sd0)))>((-(-3'sd3))?((5'sd15)<=(3'd5)):((2'd0)*(5'd11))));

  assign y0 = {3{{1{($signed(a2)>{3{p13}})}}}};
  assign y1 = (-(~(~&({p7}<<(&p12)))));
  assign y2 = (p16!=p17);
  assign y3 = (-5'sd6);
  assign y4 = (&{((p9?p5:p16)?(p10?p4:p8):(p7?p1:p10)),((&p13)?(p14?p4:p16):{p5,p2})});
  assign y5 = (((6'd2 * (p0<<b1))-((a3>a2)!=(~&p17)))>((4'd2 * {1{b2}})!=((p12>=p4)>=(a1||p5))));
  assign y6 = {{({p5,p14,p10}>={p3,p7})},(|(-{{a0,p8}})),({p17,b2,p14}<<<(+(~|p9)))};
  assign y7 = (-{2{((~&(&((p4?b1:p2))))>>>((|b2)?{p4}:{2{p6}}))}});
  assign y8 = {4{((^p14)<<<(p6>>>p2))}};
  assign y9 = (~&(~^(-2'sd1)));
  assign y10 = (+(5'd24));
  assign y11 = ((b4+p11)?$signed((a0?p9:b5)):$unsigned({1{b2}}));
  assign y12 = ((~(~(~|(5'd2 * (~&(p12<=a0))))))!=(((a2<=a1)%a3)>(&(b4<b3))));
  assign y13 = (((4'd2 * p13)<(b3))>(5'd2 * $unsigned(p1)));
  assign y14 = $unsigned((((5'd26)+(5'd10))?(6'd2 * (3'd6)):(($unsigned($unsigned((b3?p3:b1)))))));
  assign y15 = (~^p2);
  assign y16 = (~^(6'd2 * (~^(p13||p12))));
  assign y17 = ($signed(((a5/b0)<=(4'd8)))^(3'd6));
endmodule
