module expression_00878(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd2 * (4'd2))?((4'sd4)?(5'd3):(4'sd1)):((-4'sd6)!=(4'd4)));
  localparam [4:0] p1 = (~^(5'd1));
  localparam [5:0] p2 = ((-5'sd11)&&({(-2'sd1)}?{(5'd29)}:(4'sd3)));
  localparam signed [3:0] p3 = {(4'd11),(3'd4),(-4'sd4)};
  localparam signed [4:0] p4 = (5'd19);
  localparam signed [5:0] p5 = ((!(((5'd8)-(-2'sd0))<<((5'd11)<<<(2'd0))))!={4{(3'd1)}});
  localparam [3:0] p6 = (|(~^(~{(&(((5'sd6)>>(5'sd4))!=={(4'sd1),(5'sd4)}))})));
  localparam [4:0] p7 = (&(~&((-(-4'sd5))?{1{(-4'sd7)}}:{1{(-2'sd0)}})));
  localparam [5:0] p8 = (-2'sd0);
  localparam signed [3:0] p9 = (~^(-2'sd1));
  localparam signed [4:0] p10 = ((((-4'sd7)>>>(-4'sd6))%(4'd1))<=(((3'd1)===(4'd7))|(+(5'd13))));
  localparam signed [5:0] p11 = (!{2{({(4'sd2),(5'sd1),(3'sd0)}^~(-{(-4'sd0),(2'sd1)}))}});
  localparam [3:0] p12 = (4'd2 * (2'd0));
  localparam [4:0] p13 = {4{(5'sd12)}};
  localparam [5:0] p14 = {(3'sd0),(3'd6),(-4'sd4)};
  localparam signed [3:0] p15 = {(((-2'sd0)==(-4'sd0))===((5'd15)&(-2'sd0))),(((5'd0)>>>(-4'sd4))>{(3'd0)}),({(5'sd12),(5'd18)}|((4'd11)&&(5'd1)))};
  localparam signed [4:0] p16 = {(5'd4)};
  localparam signed [5:0] p17 = ({2{((3'd4)?(-5'sd14):(5'd31))}}==(((2'd1)?(4'd8):(3'd2))?((-4'sd4)<<<(2'sd0)):{4{(4'd6)}}));

  assign y0 = ({3{(-b2)}}>$signed((~|(a0<<b5))));
  assign y1 = (^{{p4,p6},$unsigned(a0)});
  assign y2 = (({((3'd2)<<(a1!=p13))})|{{(-3'sd1),(b5==b0),(4'd2 * b2)}});
  assign y3 = $signed($unsigned((+$unsigned((&{1{b1}})))));
  assign y4 = (b1?b4:b0);
  assign y5 = ({1{((p4==p10)|(p12&p6))}}!=(-{2{(p13<<p9)}}));
  assign y6 = (~&(+p17));
  assign y7 = {(&({(~&($signed((b3^~p5))))}<={(^(~&p15)),(p14?p2:b2)}))};
  assign y8 = {1{((4'd6)<(-3'sd1))}};
  assign y9 = ((b3));
  assign y10 = (~(!(~((+(|(~&p5)))||(!(p10-p0))))));
  assign y11 = (p4);
  assign y12 = {({3{b1}}&(b4?a0:b1)),{{b3,a2}},{(5'd26)}};
  assign y13 = {(~(4'd2 * $unsigned((p8&p3))))};
  assign y14 = {4{(3'd0)}};
  assign y15 = (-$signed({(5'd2 * (-(p8>=a2)))}));
  assign y16 = ((p9<<p14)%p16);
  assign y17 = ((|p11)?(~|p12):(p8?p12:p5));
endmodule
