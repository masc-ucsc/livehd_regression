module expression_00176(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|{4{(~|((2'd3)^~(4'd11)))}});
  localparam [4:0] p1 = (~|(~^(~^(~(|(4'd2 * ((4'd14)>=(4'd7))))))));
  localparam [5:0] p2 = (-3'sd3);
  localparam signed [3:0] p3 = (~^(~^(+(2'd3))));
  localparam signed [4:0] p4 = (((4'd6)+(!((3'd2)<<<(-5'sd2))))+(+((5'd7)<=(-5'sd12))));
  localparam signed [5:0] p5 = (4'd0);
  localparam [3:0] p6 = (-4'sd7);
  localparam [4:0] p7 = (-4'sd2);
  localparam [5:0] p8 = ({4{(-5'sd1)}}==(3'sd3));
  localparam signed [3:0] p9 = (((-3'sd3)?(4'd11):(-4'sd0))>={(-3'sd2)});
  localparam signed [4:0] p10 = {4{{1{{1{{2{(3'd3)}}}}}}}};
  localparam signed [5:0] p11 = ((-(~^((2'sd0)?(5'd30):(4'sd7))))?(-((4'd7)?(3'd0):(4'd8))):(|((-3'sd1)?(4'd9):(2'd3))));
  localparam [3:0] p12 = {2{{4{{1{(4'd6)}}}}}};
  localparam [4:0] p13 = {{((4'd1)?(-3'sd1):(4'd15)),((4'd15)?(4'sd7):(2'd3))},(4'd10),(2'd2)};
  localparam [5:0] p14 = ((~(-2'sd0))%(4'd10));
  localparam signed [3:0] p15 = (4'd5);
  localparam signed [4:0] p16 = ({4{((4'sd3)^~(5'd25))}}<<<({1{(2'sd1)}}?{1{(4'd10)}}:{4{(2'd1)}}));
  localparam signed [5:0] p17 = ((2'sd1)>=(|({2{(2'd1)}}==={4{(2'd2)}})));

  assign y0 = $signed({{b1,p6,a3},(+b1)});
  assign y1 = (!({3{(+b2)}}>>>(-2'sd0)));
  assign y2 = (((5'sd3)?(3'd0):{b4,p15,a5})?((2'sd0)==(p11&p9)):{1{{(2'd3)}}});
  assign y3 = ((p1>>p16)?(|{p10,p14}):(+(~|p1)));
  assign y4 = {{(~^(~^(&(!(~^a1))))),{(|{{2{p15}}})}}};
  assign y5 = {(-p12)};
  assign y6 = ({2{(2'sd1)}}<<(3'd1));
  assign y7 = $unsigned({(~&(3'sd2)),(-((b0?b5:a0)!=={a5,a2}))});
  assign y8 = (&(-((^a3)>(|p7))));
  assign y9 = (-4'sd4);
  assign y10 = (-4'sd5);
  assign y11 = ((p9>p17)%b5);
  assign y12 = ((!(-5'sd9))?((!a3)?(2'd1):(^a2)):((p12?a5:a2)<<<(3'd0)));
  assign y13 = ({3{(a0?a0:a2)}}!==(({2{b5}}?(a2<=a5):{4{a5}})^~((4'd2 * a2)?{1{a3}}:(a5?b1:a4))));
  assign y14 = (4'd15);
  assign y15 = {3{{2{{1{p12}}}}}};
  assign y16 = (((p6>>>a2))^~(a2<<b5));
  assign y17 = (({2{b1}}<(b3?p9:p16))?(3'd0):$unsigned({($signed(b4)===(a1?b0:a2))}));
endmodule
