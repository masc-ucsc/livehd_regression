module expression_00361(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~^(5'd14))||(~|(3'sd1)));
  localparam [4:0] p1 = ((((3'd6)==(5'sd12))==((3'd0)<=(2'd0)))>=(((4'd12)/(-4'sd2))>>>((5'sd5)^(-3'sd1))));
  localparam [5:0] p2 = (-4'sd2);
  localparam signed [3:0] p3 = {1{((3'd0)?(-2'sd1):(2'sd0))}};
  localparam signed [4:0] p4 = {1{((5'd24)-(-3'sd1))}};
  localparam signed [5:0] p5 = ((-5'sd1)!==(3'sd2));
  localparam [3:0] p6 = (2'd3);
  localparam [4:0] p7 = {4{(2'd3)}};
  localparam [5:0] p8 = (((3'd6)-(-2'sd1))%(4'd0));
  localparam signed [3:0] p9 = ((((-2'sd0)<(-3'sd3))==((2'sd0)>(4'd4)))<=(((4'd0)||(-2'sd0))>=((-4'sd0)==(3'd4))));
  localparam signed [4:0] p10 = {{{1{(4'd7)}},(~&(-4'sd0))},({1{(-3'sd3)}}-{(4'sd7),(3'sd1),(-4'sd2)})};
  localparam signed [5:0] p11 = (+(4'd2));
  localparam [3:0] p12 = ((&((!(5'd0))!={1{(2'sd0)}}))>>>(((-4'sd3)>>>(2'd3))&&(3'd4)));
  localparam [4:0] p13 = (^((4'd2)^(-2'sd0)));
  localparam [5:0] p14 = ((4'd4)?(3'sd2):(-2'sd0));
  localparam signed [3:0] p15 = {(((3'd3)?(-5'sd12):(5'sd12))?(|(3'd7)):((-4'sd4)?(-3'sd3):(4'sd3)))};
  localparam signed [4:0] p16 = (4'd2 * (5'd8));
  localparam signed [5:0] p17 = {2{{1{(+(~^(-3'sd1)))}}}};

  assign y0 = $unsigned({4{($unsigned(p11)>=(b1===a3))}});
  assign y1 = (5'd18);
  assign y2 = (!p0);
  assign y3 = (3'd4);
  assign y4 = (5'd2 * $unsigned((a1^b5)));
  assign y5 = ({(p17?b3:p14)}^({a1}<(a5?p6:p6)));
  assign y6 = ((((a4?a5:a3))&&$signed((a1?a2:a5)))?($unsigned(b1)?(b0<<b5):$unsigned(b2)):((p15&&a1)?(a5?b3:a4):(a4<<<a1)));
  assign y7 = (~&(5'd21));
  assign y8 = (~b2);
  assign y9 = $signed((-(~^(~&(|$signed((~^{((4'sd1)?(b4?a4:a2):(5'sd6))})))))));
  assign y10 = (4'sd6);
  assign y11 = ((!({4{(^a0)}})));
  assign y12 = (|(~^((~(~|(5'd2 * p2)))^((a4>=b4)?(~^a4):(b0<<<b4)))));
  assign y13 = ((a0===b4)?(p2&a1):{a5,a3});
  assign y14 = (p1?p10:a0);
  assign y15 = (^((-a2)?(p8?a2:a3):(3'sd1)));
  assign y16 = (~^(-5'sd5));
  assign y17 = ($unsigned(p2)?(p9):(5'sd8));
endmodule
