module expression_00609(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'sd0)&&(3'sd0))&&((4'd13)*(3'sd0)))<<<(((5'd27)<(3'd5))>=((2'd1)!=(5'd8))));
  localparam [4:0] p1 = (({((5'd24)&(-3'sd3))}!=(^((5'd4)>>>(3'd6))))&{3{{(4'd4),(-4'sd2)}}});
  localparam [5:0] p2 = {({(2'd1),(4'd8)}!==((3'sd2)&&(-3'sd1))),(((-4'sd1)<(4'd6))|{(4'sd4),(5'd25)}),(((3'sd2)!=(-4'sd0))+((-4'sd4)>=(2'd0)))};
  localparam signed [3:0] p3 = {2{{((3'd0)&&(4'd14)),{3{(-4'sd0)}}}}};
  localparam signed [4:0] p4 = (|(~&(~^{(-{(4'sd0),(-3'sd3),(2'sd1)}),((|(2'd0))!==((3'd0)?(3'd5):(3'd4))),{{(2'd0)},{(3'sd2),(5'sd9)}}})));
  localparam signed [5:0] p5 = ((-(((-2'sd0)<=(4'sd5))<<<((2'd0)&&(4'd6))))||(((5'd31)<<<(3'd6))>>((2'd3)!=(3'd0))));
  localparam [3:0] p6 = ((^((4'sd7)+(-3'sd2)))/(2'd0));
  localparam [4:0] p7 = ((5'd7)>(-3'sd0));
  localparam [5:0] p8 = ((6'd2 * ((3'd3)>=(4'd7)))+(((2'sd0)/(5'sd5))<((5'd7)%(2'd0))));
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = (-2'sd0);
  localparam signed [5:0] p11 = (-(~|((2'd0)?(-5'sd9):(4'd4))));
  localparam [3:0] p12 = (((5'sd8)?(5'd8):(4'd12))<<(5'd13));
  localparam [4:0] p13 = (3'sd1);
  localparam [5:0] p14 = (((-4'sd7)?(4'd12):(4'sd3))?((-2'sd1)<(3'd7)):{((5'd22)||(3'sd2))});
  localparam signed [3:0] p15 = {3{(3'd2)}};
  localparam signed [4:0] p16 = (+({1{((3'd0)<=((2'sd1)&(4'd12)))}}<(5'sd0)));
  localparam signed [5:0] p17 = {4{{3{(-4'sd6)}}}};

  assign y0 = (($unsigned(((a0!==a4)!={4{a0}})))!==$unsigned($signed($signed(((b4<=b4))))));
  assign y1 = ((|((~|(b2!=b2))&&({4{a3}}==(~b0))))^~((b3?a1:b0)==(5'd2 * (b0^~a2))));
  assign y2 = (+((b5?p10:b5)^(&(p7>=p0))));
  assign y3 = (a1<p15);
  assign y4 = {3{a4}};
  assign y5 = {(-5'sd10),{(|({p4,p12}<(~|p0)))},{{(2'sd1)},(&(p17>p9))}};
  assign y6 = (((p1^p3)<<(a0?p16:p10))<{4{(p2?p8:a4)}});
  assign y7 = ((^(+((a4||p15)<(p16==a3))))>=((p3^~a4)||(a3|a2)));
  assign y8 = (({4{p6}}?(b2):(p9?p12:a2))?({4{a0}}?{a3,p16,p11}:{1{p13}}):{1{$signed((a0?b1:b0))}});
  assign y9 = (~^(~({2{(~^(-b5))}}<<(~|(3'd4)))));
  assign y10 = (((b2-b2)=={4{b1}}));
  assign y11 = $signed({2{(-4'sd0)}});
  assign y12 = (3'sd2);
  assign y13 = (-4'sd3);
  assign y14 = $signed((((&(~&$unsigned(((a5?b0:b4)?(-b0):(b0>=a4))))))>(!$signed(((b1?a4:a3)?(+(b3?b1:b0)):(a2?a0:a3))))));
  assign y15 = (&(4'sd2));
  assign y16 = {3{(~a1)}};
  assign y17 = ({1{(5'd21)}}?{a2,p0}:{p13,b0,b2});
endmodule
