module expression_00997(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'sd0)<<<(-3'sd2));
  localparam [4:0] p1 = ((~&({4{(5'sd13)}}===((2'd0)==(2'd0))))!=(((2'd1)<=(3'd4))!=(&{3{(3'sd1)}})));
  localparam [5:0] p2 = {{(-3'sd2),(3'sd3),(-5'sd13)},(|{(-4'sd6)})};
  localparam signed [3:0] p3 = ({(-5'sd13),((4'd11)===(-3'sd3))}<<{((3'd7)<<<(4'd9)),{{1{(4'd8)}}}});
  localparam signed [4:0] p4 = (!(2'sd0));
  localparam signed [5:0] p5 = (-3'sd2);
  localparam [3:0] p6 = (({(3'd2),(2'sd1),(-3'sd0)}||(~&(3'd4)))-{1{(((3'd0)^~(2'd1))==((2'sd0)>=(-2'sd1)))}});
  localparam [4:0] p7 = {2{(-3'sd3)}};
  localparam [5:0] p8 = (~^(((-2'sd0)?(5'd19):(5'd24))?((2'd0)&&(5'd26)):((2'sd1)?(5'd23):(-5'sd12))));
  localparam signed [3:0] p9 = (|{3{(4'd0)}});
  localparam signed [4:0] p10 = (4'd2 * ((2'd0)<(3'd6)));
  localparam signed [5:0] p11 = (2'd3);
  localparam [3:0] p12 = {1{(((2'd1)?(2'sd1):(-3'sd2))?((3'd6)?(-4'sd3):(3'd4)):((4'd15)?(4'd5):(3'd4)))}};
  localparam [4:0] p13 = {4{((-2'sd1)^(4'd14))}};
  localparam [5:0] p14 = {(((4'd3)>>((4'sd3)!=(2'sd1)))<=(((-4'sd2)^(4'sd4))>((4'sd2)!=(3'd2))))};
  localparam signed [3:0] p15 = (2'sd0);
  localparam signed [4:0] p16 = (-3'sd0);
  localparam signed [5:0] p17 = (-3'sd3);

  assign y0 = (5'sd8);
  assign y1 = (-2'sd0);
  assign y2 = ((^(~^p3)));
  assign y3 = (5'd14);
  assign y4 = (~|((!b1)<<(&p10)));
  assign y5 = (&({p14,a0,a0}-(^(p13+p11))));
  assign y6 = ((5'sd2)|{1{((p5>=p5)!={2{p12}})}});
  assign y7 = (+(~^(&(~&({$unsigned((|(~^{(~(~(~&a1)))})))})))));
  assign y8 = (((&(4'sd6))?(-5'sd12):(b4%p13))^((5'sd1)<<(-3'sd3)));
  assign y9 = {3{((|(-3'sd3)))}};
  assign y10 = ((b4?b1:a3)^(a1!==b3));
  assign y11 = {1{{3{{2{(b4+a2)}}}}}};
  assign y12 = ((+$signed((^(a3>>a3))))!=(4'sd5));
  assign y13 = (5'd23);
  assign y14 = (^(~^(((~^b0)|{a4,a5})<(~&((a1>>a1))))));
  assign y15 = ((b2<a1)!==(a4<b2));
  assign y16 = ((2'd0)>>>(b3!=p14));
  assign y17 = (!{a1});
endmodule
