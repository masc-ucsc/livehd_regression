module expression_00028(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{({(5'sd1)}^~((4'd13)^~(3'sd3)))}};
  localparam [4:0] p1 = (4'sd6);
  localparam [5:0] p2 = (3'd0);
  localparam signed [3:0] p3 = ((-2'sd0)|(5'd8));
  localparam signed [4:0] p4 = (~|(3'd7));
  localparam signed [5:0] p5 = ((((5'sd6)==(3'sd1))&&{(4'd4),(5'd30),(-3'sd3)})?(((4'sd2)<(2'd0))===((2'd1)<<(4'sd1))):{((-5'sd13)?(2'sd1):(5'd19))});
  localparam [3:0] p6 = ((^(+(3'd2)))===(((4'd6)>>(4'd0))^(~{1{(4'd4)}})));
  localparam [4:0] p7 = (~&{4{{(5'd18)}}});
  localparam [5:0] p8 = {3{((5'd2 * (4'd8))?{2{(5'd16)}}:(2'd1))}};
  localparam signed [3:0] p9 = ({({(3'sd1),(4'd11)}<<<{(2'd1),(4'd12)})}=={3{{((-4'sd5)?(4'sd0):(4'd14))}}});
  localparam signed [4:0] p10 = ((4'd2 * ((2'd1)|(4'd10)))<=((5'sd8)-((5'd7)&&(3'sd0))));
  localparam signed [5:0] p11 = (&(~&(~&(-(~^(~|(^(~&(~&(~|(~(!(+(~^(!(3'd4))))))))))))))));
  localparam [3:0] p12 = (2'd1);
  localparam [4:0] p13 = ((((4'd0)&&(5'd15))&&((4'sd7)<<(-3'sd3)))?(-((4'd11)?(-2'sd1):(4'd14))):(((-3'sd2)&&(2'd3))^((5'd19)?(4'd9):(-2'sd0))));
  localparam [5:0] p14 = (|(~((2'd2)<=(5'd30))));
  localparam signed [3:0] p15 = ((-3'sd0)>>>(-4'sd3));
  localparam signed [4:0] p16 = (2'd0);
  localparam signed [5:0] p17 = ({3{(4'd6)}}?{((-3'sd3)?(4'sd6):(3'sd2))}:{1{(4'd2 * (4'd11))}});

  assign y0 = ({4{{4{b4}}}}!==((-(&{2{b3}}))>=((~^a2)<<{4{b1}})));
  assign y1 = (((-{2{p8}})|((p0>=p7)&&(-p3)))==(5'sd4));
  assign y2 = ((~$signed((-$signed(a1))))?(~^($signed(b1)<<(~p12))):(^(!(&(a5?b0:p2)))));
  assign y3 = (~&{2{{1{(|(-(&(+{3{b1}}))))}}}});
  assign y4 = (~^(($signed($unsigned(b0))/a1)==(~((-(^(a2-b0)))>((a1>>a3)&(a1%b2))))));
  assign y5 = (((b3/b0)>>(b3^b0))==(~(&(^b0))));
  assign y6 = $signed((~(&$signed((6'd2 * {p12,b2})))));
  assign y7 = {4{(5'sd4)}};
  assign y8 = (((p10%p6))>>((p12^p5)&(a1&&a0)));
  assign y9 = (-2'sd1);
  assign y10 = {1{$unsigned(($unsigned((5'd2 * p6))?((p1||p12)||(p11?p1:p0)):($signed(p10)|(p16&&p3))))}};
  assign y11 = (((~a4)>>(b1>=a4))===((+b5)^~{4{a0}}));
  assign y12 = ((((-2'sd0)<<(-2'sd1))-{4{p16}})|(-3'sd1));
  assign y13 = {{1{p3}},(~&a4),(a5?a5:b5)};
  assign y14 = (2'd3);
  assign y15 = (b0?p7:a0);
  assign y16 = (((!a4)?(+a3):{a1,a3,a1})?(-{(~&(~|b1))}):((|b4)&(+a4)));
  assign y17 = (4'd2 * (~(^a2)));
endmodule
