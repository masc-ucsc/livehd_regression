module expression_00659(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((!{(3'd5),(5'd21),(-4'sd3)})?(6'd2 * ((3'd7)?(2'd3):(3'd4))):(-(~&{(3'd2),(4'sd2)})));
  localparam [4:0] p1 = ((((4'sd3)<<<(2'sd1))<<(+(4'd8)))!==((-(4'd2))>=((-5'sd8)||(3'd3))));
  localparam [5:0] p2 = (((5'sd11)^~(5'd8))===(-2'sd0));
  localparam signed [3:0] p3 = (((4'sd1)&(2'sd0))<<<((3'd7)<<(5'sd15)));
  localparam signed [4:0] p4 = (&(~((~&(!(5'sd4)))<<<(|((-4'sd3)>>>(2'd0))))));
  localparam signed [5:0] p5 = {(4'sd6)};
  localparam [3:0] p6 = (~&(!(4'd8)));
  localparam [4:0] p7 = (2'sd1);
  localparam [5:0] p8 = ((~|((2'd2)?(5'sd13):(4'd11)))?{(&(-3'sd1)),((4'sd0)?(5'd4):(-5'sd4))}:{{1{{1{{2{(4'd10)}}}}}}});
  localparam signed [3:0] p9 = ((((-3'sd0)!=(3'd1))!=((5'd27)&(3'sd3)))-((~&{2{(4'd6)}})>(+(!(3'sd2)))));
  localparam signed [4:0] p10 = ({((3'd2)?(-3'sd3):(3'sd1)),{(2'd1),(4'd10),(2'd3)}}!=({((-2'sd0)>>(4'd1))}||((2'd0)?(2'sd1):(5'd6))));
  localparam signed [5:0] p11 = (~^(~^(~(3'd1))));
  localparam [3:0] p12 = (~((((2'd3)^(5'd3))<(&{2{(-5'sd12)}}))!=(|((^{1{(3'sd0)}})&&{2{(4'sd1)}}))));
  localparam [4:0] p13 = (({3{(3'sd2)}}+{(4'sd5)})<((-2'sd1)&((3'sd1)!=(4'd14))));
  localparam [5:0] p14 = ((-3'sd3)?(-3'sd0):(2'd3));
  localparam signed [3:0] p15 = ((((3'sd1)+(4'd2))|((-3'sd1)<=(4'd4)))!==(((-4'sd7)>>>(5'd26))<<((4'd15)<=(3'd4))));
  localparam signed [4:0] p16 = ((2'd2)<=(-5'sd1));
  localparam signed [5:0] p17 = (!(+(^{(^(5'd17))})));

  assign y0 = $unsigned($unsigned((-4'sd7)));
  assign y1 = ((^(&(|(3'd5))))^(&((~&(p3-p15))>{p4,p12,b2})));
  assign y2 = (b0>>a0);
  assign y3 = ($signed((^((~^a2)^~(b3))))<$unsigned(((b2%a1)*(p8^p4))));
  assign y4 = ($signed(({(p17<a0)}>>>({a3,p4})))>>((p0?p10:a4)<<$signed((b3===b0))));
  assign y5 = ({1{((-3'sd0)==={4{b5}})}}?((b5===b1)&$unsigned((a5?a3:p13))):(5'd2 * (b0?b2:b1)));
  assign y6 = (|{2{{4{(a5)}}}});
  assign y7 = (((+{3{a5}})==((~^p9)<<(a5<<<b2)))<$signed($signed((&(~&{2{(b5|b0)}})))));
  assign y8 = (((-(b3&&a1))<<((b3?b5:b1)!==(b2^a1)))===(^(5'd2 * (a2&a1))));
  assign y9 = (((b0?a3:a1)<<(a1+b1))==={3{(b2?a2:a3)}});
  assign y10 = (^{4{(p12&&p7)}});
  assign y11 = ((~&(!(a2===a2)))^{3{(&p9)}});
  assign y12 = (((p3?b5:p10)?(p17?p4:p11):(b2?p17:a2))?((p4?p15:p16)*(b3^b4)):((a3>=p14)?(p1?p3:p14):(b4?b4:p1)));
  assign y13 = ({{b2,a3},(4'd6)}?(a2?a2:a5):(b0?b3:a5));
  assign y14 = {(4'd2 * $unsigned((p8<a3)))};
  assign y15 = (&(+(5'd28)));
  assign y16 = (5'd23);
  assign y17 = (((-(~|p3))>>>(!(~p10)))?((p0?p6:p14)?(a2!=b5):(b4!==a4)):(~&((p16|p0)-(~^p4))));
endmodule
