module expression_00037(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~(-5'sd15))|(~(-4'sd5)));
  localparam [4:0] p1 = ((5'd2 * ((4'd2)|(4'd3)))|(((5'd7)?(3'd3):(2'd3))==((-4'sd4)<=(4'd13))));
  localparam [5:0] p2 = (6'd2 * (3'd6));
  localparam signed [3:0] p3 = (-3'sd2);
  localparam signed [4:0] p4 = ((-5'sd0)<<<(((-3'sd0)==(4'd1))*((3'd6)?(5'sd14):(-5'sd7))));
  localparam signed [5:0] p5 = (+{(-2'sd1),(-4'sd4)});
  localparam [3:0] p6 = ((((3'd2)?(5'sd0):(5'd10))?((2'd0)?(3'sd0):(-5'sd0)):((-3'sd3)?(4'd5):(-2'sd0)))?(((3'sd1)?(2'd2):(-5'sd10))?((4'd11)?(-2'sd0):(4'd4)):((3'd1)?(4'd2):(4'd1))):(((2'd3)?(5'd18):(-2'sd1))?((2'd3)?(-5'sd9):(5'd0)):((5'd29)?(-3'sd3):(3'sd0))));
  localparam [4:0] p7 = (5'd2 * (&((3'd7)/(4'd14))));
  localparam [5:0] p8 = ((4'd11)-((5'sd5)==(-3'sd0)));
  localparam signed [3:0] p9 = (+(-4'sd4));
  localparam signed [4:0] p10 = (+(-4'sd1));
  localparam signed [5:0] p11 = (((-2'sd1)*(2'd0))!=((-2'sd1)^~(4'd12)));
  localparam [3:0] p12 = (((5'd23)?(3'sd2):(3'd6))?(|(~|(3'd7))):(|{2{(2'd1)}}));
  localparam [4:0] p13 = {(&(~(((2'sd0)||(5'd3))&&(~&(5'd28)))))};
  localparam [5:0] p14 = {3{((2'd2)>(4'd0))}};
  localparam signed [3:0] p15 = (((-4'sd7)?(5'd14):(3'd7))>(+(2'sd1)));
  localparam signed [4:0] p16 = {((5'd26)?(2'd2):(5'd2)),((5'sd8)<=(-3'sd2))};
  localparam signed [5:0] p17 = {((2'd2)>>(-5'sd8)),{(3'd4),(2'd1)}};

  assign y0 = (-((p7||p2)*(a0!==a2)));
  assign y1 = (~(((b0>=p12)?(b0!==a0):(-p6))?(~^(5'sd11)):(~^(+(p1&&p8)))));
  assign y2 = (~(((p7>p9)?(p10?p7:p16):$unsigned((p0-p12)))&&((p8?p0:p2)&((p15)&(~|p1)))));
  assign y3 = (~^($signed((b2!==a3))<{b4,b4,b3}));
  assign y4 = ($unsigned({3{b1}})>>>{3{a0}});
  assign y5 = $signed(((&($signed((!(+$signed((^(((~b2)<<<(&a4))&($unsigned(a5)>=(+a2))))))))))));
  assign y6 = (({2{p6}}>>(~p1))<<<(~^(b4-p11)));
  assign y7 = $signed({4{((b1?a3:a3)?(p16<p17):{1{b1}})}});
  assign y8 = ((-((~&(a0<a4))-(b5*a1)))!==(+(~(&((a0>b5)+(b5|b0))))));
  assign y9 = (((p13^~p3))/a4);
  assign y10 = ((~&(p8?b4:p6))?(a0===b1):(2'sd1));
  assign y11 = ((((a4|p17)<=(b4!==a1))+(4'd2 * (p14>b0)))>>>(((b4>>p2)/b1)<<((b3-p15)%a5)));
  assign y12 = $signed($unsigned({(a2|p3),(~(~&b3)),((!b0))}));
  assign y13 = ($unsigned((((b5===b5)>>(a0^~b3))!=((a4+a1)!==(a1<<<a2))))!=(((a5&a2)>={a4})<<<($signed(b1)<<<{b3,b0,b0})));
  assign y14 = (5'd15);
  assign y15 = ($unsigned(((5'd10)?(-5'sd12):(p15>p10)))<=(&(|(-4'sd5))));
  assign y16 = (~|(|((4'd0)+(|(4'd1)))));
  assign y17 = (~|(-(4'sd2)));
endmodule
