module expression_00493(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {1{((-2'sd0)==(-3'sd0))}};
  localparam [4:0] p1 = ((((4'd1)&&(3'd7))^(~(4'd4)))^({(5'd2),(2'd0),(4'd1)}>((2'd1)>(5'd22))));
  localparam [5:0] p2 = ((6'd2 * ((4'd15)||(5'd5)))?(3'd0):(^(3'd2)));
  localparam signed [3:0] p3 = (3'd0);
  localparam signed [4:0] p4 = (2'd3);
  localparam signed [5:0] p5 = {(-4'sd0),{{(2'd3),(4'sd2)}}};
  localparam [3:0] p6 = ((((4'd12)?(4'd9):(2'd0))<<<((3'sd2)<<<(2'sd0)))?(((4'd5)-(2'sd1))*((2'd2)+(4'sd3))):(((-3'sd2)<<<(3'd3))?((4'd5)!==(2'd1)):((3'd1)?(2'd0):(3'sd0))));
  localparam [4:0] p7 = (!((4'd2 * ((2'd3)^(5'd9)))>=((2'sd1)^{(-4'sd5)})));
  localparam [5:0] p8 = (~^{(2'd2),(2'd3),(2'd0)});
  localparam signed [3:0] p9 = ((((4'sd5)!=(4'sd5))>>>((5'sd2)<(3'd7)))<<(((4'd9)^~(-5'sd3))>=((-4'sd3)===(2'd3))));
  localparam signed [4:0] p10 = ((((5'sd6)?(2'd0):(3'sd0))-((5'sd4)^(5'd7)))<=((5'd2 * (4'd14))>>>((3'd4)?(2'sd1):(3'sd1))));
  localparam signed [5:0] p11 = ((~({(3'd5),(4'd12)}+((2'sd0)?(-3'sd3):(-5'sd7))))^~(((3'sd1)?(-5'sd11):(-3'sd3))-(^(5'd22))));
  localparam [3:0] p12 = ((2'd2)&(~(-5'sd4)));
  localparam [4:0] p13 = ((((-2'sd1)?(5'd6):(4'sd4))&&((3'd2)<<(3'd1)))?{{(2'd2),(-3'sd2),(3'd6)},{(2'd0)}}:(~|({(-4'sd6),(3'd6),(3'd6)}<<((-4'sd6)>=(5'sd5)))));
  localparam [5:0] p14 = {4{(&((5'd0)^(-3'sd3)))}};
  localparam signed [3:0] p15 = (^(~(4'd15)));
  localparam signed [4:0] p16 = ({(-(4'd15)),((-5'sd1)+(2'd3))}<<(~{(4'd2),(2'sd0),(4'd13)}));
  localparam signed [5:0] p17 = ({{4{(4'd2)}},((5'd15)?(-3'sd2):(2'd1)),((2'd3)^(4'd14))}?(-3'sd3):(-4'sd2));

  assign y0 = {$unsigned({4{$signed((-a3))}})};
  assign y1 = ((6'd2 * (+(|a0)))-({(a2!==b3),(a2>>>p11)}<=(|{(p0>=b5)})));
  assign y2 = (p8!=p10);
  assign y3 = {4{a0}};
  assign y4 = (2'sd1);
  assign y5 = ((+(((b4?b5:b1)===(~|b1))>(+{3{a2}})))>(^(({3{p12}}+(-p7))<<((p15?b0:b3)|{p11}))));
  assign y6 = (p9?a2:a5);
  assign y7 = ((|(p16<b5))?(|(a1===b5)):((-a4)-(p15&p13)));
  assign y8 = $unsigned(({{{((~|b3)===(a2===b2)),$unsigned((5'd2 * a0)),{(a4),(a1&b0)}}}}));
  assign y9 = ((a2?p0:a0)!=(b3>>>a0));
  assign y10 = {3{$signed((|{1{{4{p4}}}}))}};
  assign y11 = {3{{b5,b4}}};
  assign y12 = (6'd2 * {3{p0}});
  assign y13 = (-3'sd2);
  assign y14 = {(!{(+b5),(a5<a4)})};
  assign y15 = {{1{(~^{4{b1}})}},{3{(+p3)}},{3{(a0^~b4)}}};
  assign y16 = (((a2?p14:b3)?(-a2):(-a0))?(~(&(b2?p13:p10))):((+a3)?(-a5):(^b1)));
  assign y17 = (-((!(a1?a5:p2))?((-a1)?(~a3):(~^b4)):(-(~^(~&(~|b3))))));
endmodule
