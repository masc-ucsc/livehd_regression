module expression_00808(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{(~(|(2'd1)))}}?(-3'sd1):(&(&(~&(-4'sd1)))));
  localparam [4:0] p1 = (5'sd4);
  localparam [5:0] p2 = ((-2'sd1)?(-(~(-2'sd1))):(~(-5'sd4)));
  localparam signed [3:0] p3 = {{3{{(4'd15)}}},({(4'd6),(5'd14),(5'd18)}==((5'sd0)-(4'sd3))),({3{(-5'sd12)}}<<<((4'd12)||(-2'sd0)))};
  localparam signed [4:0] p4 = (-((~&(~(-(^(^(-4'sd2))))))>((~^((-5'sd11)<<(5'd15)))<((5'd27)>=(2'd1)))));
  localparam signed [5:0] p5 = ((5'd11)-(!{(2'd3),(-5'sd0),(3'd6)}));
  localparam [3:0] p6 = (-(-(~|(~|(+(~|{3{(^(~&(4'd6)))}}))))));
  localparam [4:0] p7 = (5'd2 * (5'd22));
  localparam [5:0] p8 = ((((-5'sd9)+(-4'sd2))==((4'd15)?(4'd12):(-2'sd1)))^(((5'd7)!=(2'sd0))!==((4'd8)&(4'd1))));
  localparam signed [3:0] p9 = ((((3'd7)+(2'sd0))<={(-4'sd4),(4'sd3),(4'sd0)})>>(|(~|(3'sd1))));
  localparam signed [4:0] p10 = {1{{1{({2{((-3'sd3)>=(-2'sd1))}}&&{1{({1{(5'd18)}}<<((5'd1)>=(-5'sd10)))}})}}}};
  localparam signed [5:0] p11 = ((~^((~|(-4'sd7))||(~(3'd0))))<<<((!{4{(5'd21)}})<<<(-(~^(4'd8)))));
  localparam [3:0] p12 = {2{{2{(~|(-5'sd13))}}}};
  localparam [4:0] p13 = {((-2'sd0)^(2'sd1))};
  localparam [5:0] p14 = (~^((4'sd5)^(4'sd2)));
  localparam signed [3:0] p15 = {{3{(!(2'd3))}}};
  localparam signed [4:0] p16 = {(+(~|((-4'sd7)||(2'sd0)))),(&{(~(4'sd2))}),(((-5'sd13)>>(3'sd3))<<{(2'sd1),(4'd5)})};
  localparam signed [5:0] p17 = {3{{4{(3'd7)}}}};

  assign y0 = $signed(({{(a3!==a4)},(~^{p8,p13}),(|(p12))}^(!(6'd2 * (4'd11)))));
  assign y1 = (2'd3);
  assign y2 = (3'd6);
  assign y3 = (-3'sd3);
  assign y4 = ($unsigned((b1))>>>{b5,p11,a5});
  assign y5 = (((p6&&p2)<<<(a3|p16))>((a2^~a2)<<<(p12==a1)));
  assign y6 = (a5);
  assign y7 = (^(5'd19));
  assign y8 = (~(3'd7));
  assign y9 = (^(~b5));
  assign y10 = {4{{2{p9}}}};
  assign y11 = (5'd23);
  assign y12 = {1{{((a3!==a1)?{4{p6}}:{2{p7}}),({2{(p2+a2)}}>=({3{a3}}>>{2{p2}}))}}};
  assign y13 = (((p2?p13:a5)?(p2>b3):(b5|b3))-(6'd2 * (a1>>p12)));
  assign y14 = ((!{4{a0}})?{2{{3{a3}}}}:{3{(-p10)}});
  assign y15 = (~^((!(-2'sd0))!==((-3'sd2)<((~^a4)-(a5==b4)))));
  assign y16 = (3'sd2);
  assign y17 = (((p8|p11)+(+p11))<=((p0||p8)^{a1,p5}));
endmodule
