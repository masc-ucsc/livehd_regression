module expression_00227(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd0);
  localparam [4:0] p1 = {(((3'd1)===(3'sd2))^~((4'd15)==(5'd11))),(4'd5)};
  localparam [5:0] p2 = ((-4'sd6)>>(-4'sd5));
  localparam signed [3:0] p3 = (((4'd1)!==(3'd4))*((5'd15)|(3'sd2)));
  localparam signed [4:0] p4 = (4'd11);
  localparam signed [5:0] p5 = (4'd6);
  localparam [3:0] p6 = ((+((|(-5'sd0))&&((2'd0)&(3'd5))))>>>(^(((2'd3)/(-5'sd14))<=(5'd2 * (5'd30)))));
  localparam [4:0] p7 = (-{2{(-(^(&{3{(3'd7)}})))}});
  localparam [5:0] p8 = {3{(^((~&(3'd2))<={3{(5'd17)}}))}};
  localparam signed [3:0] p9 = (4'sd7);
  localparam signed [4:0] p10 = {2{(-4'sd5)}};
  localparam signed [5:0] p11 = (4'sd1);
  localparam [3:0] p12 = (+((|(-(((3'd4)?(5'sd0):(4'd15))?((5'sd5)?(5'sd3):(4'sd4)):((5'sd10)|(-5'sd10)))))<((&((4'd11)?(5'd10):(3'd4)))^~((3'd0)?(4'd10):(4'd13)))));
  localparam [4:0] p13 = (((2'd1)<=(3'd4))>=(~|(3'd7)));
  localparam [5:0] p14 = {(4'd4),(5'd9),(4'd2)};
  localparam signed [3:0] p15 = ((5'd18)?(5'd2):(4'd11));
  localparam signed [4:0] p16 = (~(((-2'sd1)?(4'd1):(2'sd0))?(4'd13):((3'sd0)?(-2'sd0):(5'd9))));
  localparam signed [5:0] p17 = ({{(2'd3)},((3'd2)>=(2'd3))}!=={{(-4'sd3),(5'd27),(-4'sd3)},((5'd17)?(5'd18):(2'd0))});

  assign y0 = (~|(2'sd0));
  assign y1 = {((p0+p0)>>>{p9,p6}),({p10,p5,p11}?(p4==p11):(p10^p13))};
  assign y2 = (-4'sd3);
  assign y3 = (^((2'sd0)&&(-2'sd1)));
  assign y4 = (5'd12);
  assign y5 = (5'd24);
  assign y6 = {2{(+(4'd12))}};
  assign y7 = ((|b3)!=(^a2));
  assign y8 = (4'sd4);
  assign y9 = (p3==p1);
  assign y10 = ({1{{a5,p17,b5}}}!=(b3?a0:a5));
  assign y11 = $signed(((p1<<p0)?((p5?p14:p5)):(~(p0))));
  assign y12 = ((-4'sd6)+(p1<<<p3));
  assign y13 = ({(p3?p17:p10),(p5!=b0)}<=(^(((a5)!==(a2)))));
  assign y14 = {((a1!==b0)!==(5'd2 * a1)),((!p2)>=(a2<p15)),{(&a1),(+b4),(b0-a1)}};
  assign y15 = {3{{4{{3{b5}}}}}};
  assign y16 = ((-($signed((-{3{p9}}))?((^(+a0))===(b3?b0:a5)):{{p5,p7,p8},{1{(~^p7)}}})));
  assign y17 = ((|((a2!=a4)|$unsigned(a1))));
endmodule
