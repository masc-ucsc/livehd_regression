module expression_00638(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'sd1)?(4'sd4):(-3'sd2))?{1{(2'd2)}}:((-2'sd1)?(2'sd1):(5'd15)))?{3{((5'd31)+(2'd3))}}:(((3'd5)?(2'sd1):(5'sd7))?((5'd4)?(4'd7):(3'd6)):((2'sd0)?(4'd13):(5'sd0))));
  localparam [4:0] p1 = (((!(2'd0))>>((4'd10)&&(5'd19)))-{3{(4'd9)}});
  localparam [5:0] p2 = ((((2'd1)&&(5'sd9))<<<{(4'd10),(5'd21),(-5'sd0)})|(((2'd1)?(5'sd12):(5'd20))?((3'd7)<<<(-2'sd1)):{(-5'sd15)}));
  localparam signed [3:0] p3 = (5'sd6);
  localparam signed [4:0] p4 = (((3'sd1)?((4'd7)?(5'd26):(2'sd1)):(-(5'd18)))==((2'd3)!=(-3'sd3)));
  localparam signed [5:0] p5 = (4'd12);
  localparam [3:0] p6 = ((2'sd1)<<{((3'sd3)|(-4'sd2)),((5'd17)>(-3'sd0)),((-3'sd1)!==(5'd18))});
  localparam [4:0] p7 = ((3'd6)-(5'd29));
  localparam [5:0] p8 = {4{(-3'sd2)}};
  localparam signed [3:0] p9 = (2'sd0);
  localparam signed [4:0] p10 = ({1{(-5'sd11)}}<=((3'd5)+(4'sd3)));
  localparam signed [5:0] p11 = ((((2'sd0)-(2'd2))^~((-4'sd4)+(-5'sd9)))<<((2'sd0)|((2'd3)+(4'd1))));
  localparam [3:0] p12 = (~&(((5'sd12)?(5'd12):(-3'sd1))>>(^(~|(2'sd1)))));
  localparam [4:0] p13 = (-(+(^(~^(~^((^((3'sd2)|(4'sd2)))!==(((-5'sd13)<(-4'sd0))||((2'd2)==(2'sd1)))))))));
  localparam [5:0] p14 = (5'sd9);
  localparam signed [3:0] p15 = ({2{(2'sd1)}}?((4'sd6)?(2'd2):(2'd2)):{3{(2'd2)}});
  localparam signed [4:0] p16 = {1{(~|(|{({{1{(-4'sd1)}}}|((4'd7)?(5'd3):(5'sd4))),(+((~|(3'd1))?{3{(3'd4)}}:((3'd0)?(4'd10):(2'sd1))))}))}};
  localparam signed [5:0] p17 = (~(3'd4));

  assign y0 = {4{(~&a0)}};
  assign y1 = (~|(((^(p11?a0:p6))?(!$signed(b5)):(p16-b4))>>>(&(-((p15^~b5)?$unsigned(p17):(&a3))))));
  assign y2 = {((~&(|((+a1)>>>(b4|a3))))),{(!(6'd2 * (!(p2>=p6))))}};
  assign y3 = ((^((+(~&p11))!=(|{p2,p2,p7})))+(!((2'sd0)+(~|(b5<<<p6)))));
  assign y4 = (((2'd0)>>(a1===a1))?((-3'sd1)?(p8^~p1):(-5'sd13)):((-2'sd0)<<(p13-p2)));
  assign y5 = {3{{2{(p4+b5)}}}};
  assign y6 = (4'd8);
  assign y7 = (^(~|(p17^~b1)));
  assign y8 = (p17==p17);
  assign y9 = (((~^(b0<<a2))&&((a3?a5:a1)>=(a5>>b1)))<(~((~&(b3?b0:b0))-(b3?a2:b2))));
  assign y10 = (((b2<=p13)?(p4||p16):(b1?p14:a2))?((!(a0>>>p10))<<(b5?p11:b5)):(+(5'sd13)));
  assign y11 = {2{({(4'd7)}^~{3{b2}})}};
  assign y12 = (|(((!$signed(b3))>>>(~{p2,a3}))<(!(~&(3'd2)))));
  assign y13 = (((-4'sd0)?$signed((p5>=p4)):(p7?p7:p14)));
  assign y14 = (3'd3);
  assign y15 = (-2'sd1);
  assign y16 = (({1{(({(~^a4)}>>(a0<<p15)))}}));
  assign y17 = $signed((((b3?p16:b2)?$unsigned(a5):$signed(a4))^~((a0?a4:a4)?$signed(a0):$signed(b5))));
endmodule
