module expression_00919(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&{2{((-5'sd3)===(5'sd2))}});
  localparam [4:0] p1 = ((-(|{((3'sd1)<<(-2'sd0))}))^~{{(~^(!(~(-4'sd7))))}});
  localparam [5:0] p2 = ((((3'd0)?(-4'sd7):(5'sd5))>=((5'd2)!=(-3'sd3)))===(((5'sd10)!=(5'sd7))?((-4'sd7)>(-4'sd4)):((5'sd2)<<<(-3'sd0))));
  localparam signed [3:0] p3 = (~^(2'd2));
  localparam signed [4:0] p4 = {{{(2'sd0)},{(-3'sd2)},{(2'd3),(3'd1)}},{{{(-5'sd15),(-3'sd2),(-4'sd1)},{(-2'sd0)}}},{{{(3'd7),(5'd7),(3'sd0)}}}};
  localparam signed [5:0] p5 = ((&{4{((4'd2)!=(5'd28))}})>>(((3'd0)&&(2'sd1))^((5'sd14)>(3'sd3))));
  localparam [3:0] p6 = (2'sd1);
  localparam [4:0] p7 = {4{(4'd7)}};
  localparam [5:0] p8 = ((~(~^(+(-{((4'd2)<<<(4'sd6)),((2'd2)<(-3'sd2))}))))+((-(&{(-5'sd12),(3'd3),(4'd10)}))<<<(((-4'sd5)<<<(-5'sd10))^(~^(5'd13)))));
  localparam signed [3:0] p9 = {1{(((5'd29)?(2'sd1):(5'sd9))?((-3'sd0)&(2'sd1)):(5'd2))}};
  localparam signed [4:0] p10 = ({4{(4'd5)}}?(~^(2'd0)):((4'd15)?(4'sd3):(4'd13)));
  localparam signed [5:0] p11 = ((3'd5)>>(-4'sd6));
  localparam [3:0] p12 = (-3'sd2);
  localparam [4:0] p13 = ((2'd0)?(2'sd1):(5'sd4));
  localparam [5:0] p14 = {1{(6'd2 * ((5'd17)^~(3'd5)))}};
  localparam signed [3:0] p15 = ((((3'd6)<(4'd15))?{3{(5'sd8)}}:((4'sd2)?(2'sd1):(-2'sd1)))>={((5'sd5)?(-4'sd3):(-2'sd1)),((2'd1)<=(4'd14))});
  localparam signed [4:0] p16 = (((|(3'd5))?((-2'sd0)&(3'sd1)):((3'sd2)<<<(5'd21)))?(((2'd1)>>(-3'sd2))>={(4'd2),(4'd15),(5'd2)}):((~|(4'd1))<<<((3'd6)>>>(3'd0))));
  localparam signed [5:0] p17 = (!{2{((&(-5'sd11))?{4{(2'd0)}}:(&(-2'sd1)))}});

  assign y0 = ((((~&p5)%a0)||((b3>>a4)<(b3&&b4)))==(((!a1)/a5)<((a1>=a4)<=(p8-b2))));
  assign y1 = ((!(5'd17))?(+(&(~^(!(p15?b0:a4))))):$unsigned(((5'sd15)?(-3'sd3):(3'sd2))));
  assign y2 = {{(((5'd9)&&{(b1-p16),(p1<=b0)})>>(2'd1))}};
  assign y3 = {(b4),(p5?b2:p16),(p11?p0:p4)};
  assign y4 = ((^$signed($signed(a1)))<<<(|$signed((b0?b1:b5))));
  assign y5 = (($signed($signed($unsigned(p15)))^(b0?a3:b2))>>$signed($signed(((b1*b2)<=(b2===b2)))));
  assign y6 = (({2{b4}}?(a5<<a0):(a2<<<p9))?{2{(a1-b3)}}:((5'd2 * b0)===(!a5)));
  assign y7 = (4'd10);
  assign y8 = (~|((3'd0)>>>$unsigned({(|{p15})})));
  assign y9 = (-(3'sd2));
  assign y10 = (((a4?a1:a3)&&{a2,b0})!==(|(~|{{(b3?b3:b2)}})));
  assign y11 = {4{({1{p8}}==(p3))}};
  assign y12 = ((~$unsigned((^b0)))==({2{a5}}<=(b0!=a0)));
  assign y13 = {4{p17}};
  assign y14 = (~|{2{((&(~&(!p2)))^~({4{p13}}!=(p16>>>p13)))}});
  assign y15 = (~|($unsigned({b1,b2})?$signed((p0<b3)):(+(b5!=b3))));
  assign y16 = (+(p15^~a0));
  assign y17 = ((+(b1?p9:p2))?(-2'sd1):((^a1)===(a5>a5)));
endmodule
