module expression_00428(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(-4'sd3)}};
  localparam [4:0] p1 = (5'd0);
  localparam [5:0] p2 = ((~&(2'd3))!==(5'd0));
  localparam signed [3:0] p3 = ((((3'd0)?(5'sd11):(5'd25))>(-3'sd3))?(4'd11):(|{(~|(3'sd2))}));
  localparam signed [4:0] p4 = (&(+(&{{(|(-2'sd1)),(~&(2'd3))}})));
  localparam signed [5:0] p5 = (((-3'sd3)<=(-2'sd0))>>>(((3'd0)==(5'd4))-(-2'sd1)));
  localparam [3:0] p6 = (((|(3'sd2))?((4'd4)>>(4'd6)):(~&(2'd3)))&(((5'sd10)<=(3'd6))==((4'sd6)>(3'sd3))));
  localparam [4:0] p7 = ((((4'sd2)^~(3'd2))>((5'sd1)|(3'd1)))>(((3'd6)!=(2'd3))===(-(&(2'd0)))));
  localparam [5:0] p8 = ((((5'sd1)/(4'd9))>>((5'd16)>(-4'sd5)))|(((3'd7)!=(5'd9))!=((3'd1)%(3'sd3))));
  localparam signed [3:0] p9 = (6'd2 * ((3'd7)<<(2'd1)));
  localparam signed [4:0] p10 = {(~((4'd3)>(4'd8))),(2'd2)};
  localparam signed [5:0] p11 = {4{(5'd5)}};
  localparam [3:0] p12 = {1{(~(~&(3'd3)))}};
  localparam [4:0] p13 = (-4'sd2);
  localparam [5:0] p14 = {2{(4'd7)}};
  localparam signed [3:0] p15 = {((^{(4'sd5)})-{(2'd3),(3'd1),(2'd1)})};
  localparam signed [4:0] p16 = ((((3'd2)<=(4'd10))|{1{(2'd1)}})>>>((~^(-4'sd5))!=((4'd5)!=(-4'sd1))));
  localparam signed [5:0] p17 = ((((2'sd1)+(-2'sd1))<<<(3'd1))>>>(5'd12));

  assign y0 = (~&{3{{(-b4),(|b1),(!p14)}}});
  assign y1 = {{(p4?p13:p6)}};
  assign y2 = {4{p8}};
  assign y3 = {{{(&p13),(p0<<p3),(-p0)}}};
  assign y4 = ({({{p4,p2,b4}}-(p3==p13))}^({(p13<p7),(b1<=p16)}>((b0-a5)>={p7,p11,p9})));
  assign y5 = (^(~(~&((-(p5^~p10))&&(+{p0,p17})))));
  assign y6 = {4{{(&{{3{b4}}})}}};
  assign y7 = $unsigned({1{((((p0|p9)?(p10^p17):(4'd2 * p8))||{3{{4{p0}}}}))}});
  assign y8 = {(({p1}<<(p13>>p0))<<((~p1)=={p13})),(({p17,p5,p3}<=(p17&&p16))&&({p5,b1,p2}&&(~|p3)))};
  assign y9 = (((p1&&p16)?{3{p12}}:(~&p6))>(4'd13));
  assign y10 = $unsigned(p1);
  assign y11 = ((~|b2)&&(!p10));
  assign y12 = (((p3&p17)<<<{1{(p0?p15:p15)}})<=({1{(-3'sd2)}}&{1{(p8>>p6)}}));
  assign y13 = (+(~|(|(p13?p2:p17))));
  assign y14 = (~(|(({p8,a3})>=(^(b3!=a2)))));
  assign y15 = (!(2'sd1));
  assign y16 = (2'd0);
  assign y17 = $signed((({(3'sd2),(-2'sd1),{b5,a1}}<=(!((-3'sd1)&&(p6))))));
endmodule
