module expression_00749(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{{(4'd5),(4'sd3),(-3'sd1)}}}<=((-4'sd4)?(2'sd1):(2'd2)));
  localparam [4:0] p1 = (-(!(-5'sd3)));
  localparam [5:0] p2 = {{3{(3'sd3)}}};
  localparam signed [3:0] p3 = {{{(2'd1),(2'sd0)}},{((2'd3)?(5'd20):(2'd3)),((2'sd0)?(-3'sd2):(-5'sd5))},(((-5'sd9)==(4'd1))&&((5'd21)?(3'sd3):(5'sd14)))};
  localparam signed [4:0] p4 = ({2{(~^(+(4'd3)))}}==(!{4{((-2'sd1)<<(4'd15))}}));
  localparam signed [5:0] p5 = (~|{(-5'sd9),(2'd1)});
  localparam [3:0] p6 = {(~|(5'd27))};
  localparam [4:0] p7 = {(~^({(2'd1),(2'd0)}<<<(3'd2))),(2'd0)};
  localparam [5:0] p8 = ((2'd0)^~(4'd0));
  localparam signed [3:0] p9 = ((6'd2 * ((2'd2)?(3'd6):(2'd1)))>>{(2'd1),(^(3'sd2)),((4'sd4)>>>(2'd2))});
  localparam signed [4:0] p10 = (((5'd8)&(3'd1))?(!(|(2'sd1))):((5'd9)?(3'd1):(-3'sd1)));
  localparam signed [5:0] p11 = (!((+(~&(-((2'd0)^(4'sd1)))))>>>(((-2'sd1)>>(3'd5))^(&(5'd26)))));
  localparam [3:0] p12 = (~^{2{(|(~&((~^(3'sd1))+(+(2'sd0)))))}});
  localparam [4:0] p13 = {1{{4{{2{(3'd2)}}}}}};
  localparam [5:0] p14 = (((-3'sd0)<=((3'sd1)+(2'sd0)))?(3'sd1):(((3'd0)===(5'd1))||((5'd22)>=(3'd2))));
  localparam signed [3:0] p15 = (4'd2 * {(3'd0),(2'd3),(2'd0)});
  localparam signed [4:0] p16 = {(!{(2'sd1),(3'd7),(3'd0)}),(~&((2'd1)?(3'd1):(-2'sd0))),{2{(-5'sd6)}}};
  localparam signed [5:0] p17 = (2'd3);

  assign y0 = (4'd8);
  assign y1 = {{3{(b5<<a2)}}};
  assign y2 = (((b3?p8:a5)/a2)<<(b3?a1:p13));
  assign y3 = ((3'd0)>>>(b5>>p1));
  assign y4 = ((b0-p10)&&(a1>>a5));
  assign y5 = (|(~&((~^(~|b3))&(4'sd7))));
  assign y6 = (2'sd1);
  assign y7 = (5'd2);
  assign y8 = $signed({(p17|a0)});
  assign y9 = ($signed(((p17+p8)&&(a2==a1)))^~$unsigned($unsigned((((p17))&($signed(p9))))));
  assign y10 = (4'd6);
  assign y11 = {{{(a0!==b0)},(~(&p0))},(!(~&((b1>=p6)!={b5})))};
  assign y12 = (~(~|(((p10?p14:p8)==$signed({2{p14}}))&((p8?p7:p8)<<$signed((+{2{p17}}))))));
  assign y13 = (4'd2 * (a0===a2));
  assign y14 = (5'd15);
  assign y15 = {b2};
  assign y16 = (~(~|(((5'd2 * (a2<<<a0))&((^b5)<<(5'd2 * a1)))||(((~&b5)<(b4+b2))>=((b1^~b4)<=(a2!=a1))))));
  assign y17 = {$signed({{2{a3}},(p16<<a2),{1{(b3?a1:p5)}}}),{4{(!(b0))}}};
endmodule
