module expression_00804(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~&((3'sd1)?(-5'sd14):(4'd9)))?((-(-3'sd0))?(~|(-2'sd1)):((5'd12)?(3'd0):(4'sd2))):(~(~|((3'd6)?(4'd6):(-2'sd1)))));
  localparam [4:0] p1 = ((2'd2)?(^((-4'sd0)|(5'sd5))):(6'd2 * (4'd14)));
  localparam [5:0] p2 = (!((~|(!(|((3'd2)>(3'd5)))))&(((2'sd0)>>(2'd2))*(|(3'd1)))));
  localparam signed [3:0] p3 = ((((-4'sd3)?(2'd0):(-2'sd1))<=(4'd10))==(((4'd14)?(3'sd1):(5'd6))?((-4'sd0)?(5'sd14):(4'sd6)):((2'd1)/(4'd7))));
  localparam signed [4:0] p4 = (((5'sd8)?(3'sd3):(3'd5))?{2{(5'd8)}}:{3{(-4'sd3)}});
  localparam signed [5:0] p5 = (((2'sd1)?(2'sd1):(4'd4))===(((4'sd0)||(-3'sd0))>((4'sd4)+(5'd13))));
  localparam [3:0] p6 = (((5'd26)-(4'd5))+((2'sd0)<=(5'sd10)));
  localparam [4:0] p7 = (-{{{(3'sd3)}},((5'd9)>>>(-4'sd0))});
  localparam [5:0] p8 = ({(!((5'd4)-(5'd29)))}&(~&(|((3'd1)&&(4'sd3)))));
  localparam signed [3:0] p9 = (^(2'd2));
  localparam signed [4:0] p10 = ((4'd10)&(4'd2 * (2'd1)));
  localparam signed [5:0] p11 = {(5'd4)};
  localparam [3:0] p12 = ((~&((-4'sd3)!==(5'd9)))===(~{2{(5'sd0)}}));
  localparam [4:0] p13 = (((-2'sd0)?{(-3'sd3),(5'd4),(3'd5)}:((3'd7)?(2'd2):(2'd0)))>{2{{2{(5'sd7)}}}});
  localparam [5:0] p14 = ({3{(2'sd0)}}==((4'd13)==={1{((-4'sd6)?(-5'sd5):(5'd21))}}));
  localparam signed [3:0] p15 = (((-5'sd13)?(2'sd1):(-3'sd2))?((-4'sd7)?(2'd3):(2'd0)):{(-3'sd3)});
  localparam signed [4:0] p16 = (~(&((4'd14)?(3'd0):(-3'sd1))));
  localparam signed [5:0] p17 = (((-3'sd2)+(5'd29))/(2'd1));

  assign y0 = (~(5'd7));
  assign y1 = (({2{(p9&&p4)}}<{4{a4}})>{3{{1{(p4<=a3)}}}});
  assign y2 = {{2{(p0&p3)}}};
  assign y3 = (4'sd5);
  assign y4 = (a5^~a3);
  assign y5 = ({1{({2{(p8<<b1)}}+(b5?p8:a1))}}^~(((p1?b3:p17)||(p15+a3))<=((p16?b5:a5)>(p9>>>a4))));
  assign y6 = {3{{2{(a2!==a2)}}}};
  assign y7 = (2'd1);
  assign y8 = (~|({({p12,p9,b5}?(a2?b2:a5):{b5,b4,a2})}?(~|(~^((a4?a4:a1)?(b4?b3:a3):{a3}))):({b3,p5,a3}?{a3}:(^a0))));
  assign y9 = ($signed((((b0>>a4)<=(a5^a1))))<<(((b4!=a1)<=(a5===b1))));
  assign y10 = ((~^(-((p2>=b0)|(~|p2))))^((~(-p1))&(a5&&b5)));
  assign y11 = (!{2{{2{(-(a1?a3:b5))}}}});
  assign y12 = (4'sd6);
  assign y13 = {2{b1}};
  assign y14 = (5'd10);
  assign y15 = (~&(p2&b2));
  assign y16 = ({3{$signed(a5)}});
  assign y17 = ((-4'sd2)<<<((b1)===(-5'sd0)));
endmodule
