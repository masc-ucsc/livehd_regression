module expression_00903(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd5)/(-2'sd0))||(~((-5'sd8)>(-3'sd2))))&&(~^(|(~|((~&(-2'sd0))<<<(^(4'sd2)))))));
  localparam [4:0] p1 = (~(~^((((2'd0)^~(-3'sd3))^((5'd26)>(5'd12)))&{4{{(4'd2)}}})));
  localparam [5:0] p2 = (((4'd6)?(3'd3):(4'd12))?((2'd3)?(4'd11):(2'sd1)):((3'sd1)?(2'sd0):(-5'sd6)));
  localparam signed [3:0] p3 = ((3'sd1)>>>(4'd13));
  localparam signed [4:0] p4 = (5'd2 * ((5'd7)&&(5'd14)));
  localparam signed [5:0] p5 = (-((((-3'sd3)?(-5'sd5):(-3'sd2))&(5'd8))?{((2'd1)!=(-4'sd5)),((5'd2)-(3'sd0))}:{((2'd2)?(-2'sd1):(2'd3)),((3'sd1)?(4'd13):(5'd20))}));
  localparam [3:0] p6 = {(5'sd12),(~(2'sd0))};
  localparam [4:0] p7 = (-((&(~((3'd4)?(2'd1):(-2'sd1))))?{{{(3'd2),(5'd3)}}}:{1{(-(|{2{(3'd7)}}))}}));
  localparam [5:0] p8 = {(3'sd0)};
  localparam signed [3:0] p9 = ((~^{(2'sd1),(3'd4),(3'd2)})^~{(-3'sd1),(4'd9)});
  localparam signed [4:0] p10 = ((((4'sd1)>>(5'd15))!==(^(|(-2'sd1))))&&(((4'd3)<=(-3'sd1))^~((2'd2)^~(-2'sd0))));
  localparam signed [5:0] p11 = (3'sd2);
  localparam [3:0] p12 = ((((5'sd6)>>>(2'd2))||((3'd7)==(5'd3)))===(((4'd0)+(-4'sd2))*((5'sd7)===(-2'sd1))));
  localparam [4:0] p13 = (3'd3);
  localparam [5:0] p14 = {4{{1{(-2'sd1)}}}};
  localparam signed [3:0] p15 = {4{((3'sd2)||(4'sd1))}};
  localparam signed [4:0] p16 = (~^(&{{(4'sd1),(-3'sd0),(2'd3)}}));
  localparam signed [5:0] p17 = (!(&(~^(-2'sd0))));

  assign y0 = ((~(a4===b3))<((p2==p5)==(p8>p15)));
  assign y1 = (-3'sd3);
  assign y2 = ((-({4{p15}}-(&(3'd2))))>>((b4===b1)-(p16>=a2)));
  assign y3 = {{1{(4'd2)}},(4'd11)};
  assign y4 = {(5'd4)};
  assign y5 = (~^(~{2{({3{p14}}||{4{a5}})}}));
  assign y6 = (2'd3);
  assign y7 = ({{(p16!=a1),{p16,p5,a3},{a1,a5}},({b3}^~(b3|p17))}>{(((p0!=a4)^(b4<<p17))|({a2}^~(p7||a5)))});
  assign y8 = ((~|(~^b1))==(b1<=b4));
  assign y9 = (((~^(a3^~b4))%b3)<((~^((a4&b4)>>(b5<=p16)))&((a1>>b1)/p3)));
  assign y10 = $unsigned((((~&(a1?a0:a0))!==$unsigned($signed($signed((a3)))))^~$signed((-(($signed(p3)^(6'd2 * p8))>=((p2<<p0)>(p1^p2)))))));
  assign y11 = (-5'sd14);
  assign y12 = (-3'sd0);
  assign y13 = (-2'sd0);
  assign y14 = (3'd7);
  assign y15 = ($unsigned(a1)?(&b4):(4'd0));
  assign y16 = {((a2==a0)<<<{a4}),(b2?a0:a5)};
  assign y17 = {(&(a1-p9)),(+(-4'sd5))};
endmodule
