module expression_00504(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(+({(4'sd4),(2'd3)}!=(^(5'd19)))));
  localparam [4:0] p1 = (-4'sd3);
  localparam [5:0] p2 = {3{(3'sd2)}};
  localparam signed [3:0] p3 = {(4'd7),((3'sd0)>=(2'd1))};
  localparam signed [4:0] p4 = (((2'd1)^~(3'sd1))?((2'd0)/(-2'sd0)):((2'd0)&&(5'd23)));
  localparam signed [5:0] p5 = {2{(((-5'sd13)!=(5'd3))+{4{(5'd26)}})}};
  localparam [3:0] p6 = {(5'sd2),{(3'd3),(-5'sd15),(2'd2)},(4'd15)};
  localparam [4:0] p7 = {4{{4{(3'd7)}}}};
  localparam [5:0] p8 = (~^((((3'd7)?(3'sd0):(4'sd1))?((5'd28)>>>(4'd5)):((5'd2)^~(-5'sd2)))<(((3'd6)?(2'd0):(3'd7))>>((3'sd3)<<(4'sd2)))));
  localparam signed [3:0] p9 = (-(2'd3));
  localparam signed [4:0] p10 = {1{({4{(^(4'sd7))}}===({1{(~&(5'd0))}}&&(^{1{(4'sd0)}})))}};
  localparam signed [5:0] p11 = (2'd2);
  localparam [3:0] p12 = (-{(5'd0),(-3'sd3),(2'sd0)});
  localparam [4:0] p13 = (((-2'sd1)?(-4'sd3):(-5'sd7))?(((2'sd0)?(2'sd1):(4'd6))^((4'sd7)===(4'd9))):(((-2'sd1)===(-5'sd1))-((-4'sd0)?(-5'sd10):(5'd20))));
  localparam [5:0] p14 = (((4'd0)?(-2'sd1):(3'd7))?(((3'sd0)^(2'sd0))&&((5'd7)&(2'd3))):((4'd6)-(5'd2 * (4'd11))));
  localparam signed [3:0] p15 = {2{{3{((2'sd0)^~(3'd1))}}}};
  localparam signed [4:0] p16 = (+(+(2'sd0)));
  localparam signed [5:0] p17 = {{1{({2{(4'd13)}}>>>{1{(-4'sd0)}})}},(3'd7),{{((3'd3)!==(2'd3)),{3{(4'd15)}}}}};

  assign y0 = {1{(5'd19)}};
  assign y1 = ((b2&a3)%p13);
  assign y2 = (|b0);
  assign y3 = $unsigned((5'sd9));
  assign y4 = ((|$unsigned((6'd2 * (5'd31))))^~{{{p7,p0,p10},($unsigned(p16)),(5'd28)}});
  assign y5 = (5'd20);
  assign y6 = {1{((((p15?p13:p6)^{3{p12}})!={2{{1{p3}}}})^~{1{({1{(a1?b0:a5)}}===(a3?b2:b1))}})}};
  assign y7 = {1{$signed((($signed(((4'd2 * b1)))<=(~|(~&{2{b4}})))))}};
  assign y8 = ((p17%a2)?(a1%a3):(p0|b5));
  assign y9 = {1{(~(~^(({2{(&$signed((~|({2{p10}}?{1{p17}}:{3{p17}}))))}}))))}};
  assign y10 = (~|(|(+{2{{(p9<<b1)}}})));
  assign y11 = {{p11,b4,a0},(a0<=b2),(3'd1)};
  assign y12 = (|((~{2{{a5}}})));
  assign y13 = $signed($signed($signed((2'd3))));
  assign y14 = ((|(+(|((^{3{p11}})^(a5-p15)))))^(|((!(p0>>b1))&(+(b1===b3)))));
  assign y15 = (-($signed({4{(~^a2)}})+(-{4{(p6<=p17)}})));
  assign y16 = {2{(({a2}===(a1>=a5))>={(|p3),(~^p11)})}};
  assign y17 = ((5'sd8)>=(p13!=a1));
endmodule
