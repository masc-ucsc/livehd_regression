module expression_00970(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd2 * (2'd3));
  localparam [4:0] p1 = ((((4'sd2)?(2'sd0):(-4'sd6))<<<((2'sd1)?(-3'sd2):(5'd29)))>>((((-2'sd0)?(4'd15):(3'sd1))-((3'd2)>>(3'sd1)))!==((-3'sd3)?(5'sd1):(5'd2))));
  localparam [5:0] p2 = (4'sd5);
  localparam signed [3:0] p3 = ((2'd2)?(3'd7):(-5'sd7));
  localparam signed [4:0] p4 = (~^(4'sd1));
  localparam signed [5:0] p5 = ((-5'sd9)>>((~(4'sd1))<=((5'sd7)+(5'd24))));
  localparam [3:0] p6 = ((((3'd4)|(4'd12))<<((5'sd8)<<<(5'd14)))<<<(((-3'sd0)|(5'd10))>>((2'd0)<(2'd1))));
  localparam [4:0] p7 = (-5'sd2);
  localparam [5:0] p8 = (+(((2'sd1)|((2'sd1)?(2'd1):(3'd6)))-(((5'd18)<=(2'd2))?((3'sd2)>>>(2'd1)):(&(-3'sd2)))));
  localparam signed [3:0] p9 = {2{(-5'sd2)}};
  localparam signed [4:0] p10 = {4{(3'sd0)}};
  localparam signed [5:0] p11 = (((5'd21)<(2'd1))&&((-2'sd1)^~(5'sd3)));
  localparam [3:0] p12 = ((((3'd5)!=(4'd12))?((2'd2)^(-2'sd0)):((3'd6)>>>(2'd2)))?(((5'sd10)?(-2'sd0):(-2'sd1))?((-5'sd3)+(4'd12)):((3'd0)?(-2'sd0):(2'd0))):(((2'd2)*(4'd1))===((-3'sd3)*(2'sd1))));
  localparam [4:0] p13 = ((-2'sd1)!=((4'd14)^((3'd7)>=(2'd0))));
  localparam [5:0] p14 = ((-3'sd0)?(4'sd6):(3'd0));
  localparam signed [3:0] p15 = (~|(((4'd2)?(5'd21):(-2'sd0))?(~(5'sd11)):((5'sd0)?(-2'sd0):(2'd3))));
  localparam signed [4:0] p16 = (&{4{(+{1{{3{(3'd4)}}}})}});
  localparam signed [5:0] p17 = (+((&(5'd17))<<<((2'd1)>>>(4'd5))));

  assign y0 = (|({((&(p11))),((b4?p5:b4))}));
  assign y1 = ((~^(!(~|(3'd5))))<(3'sd2));
  assign y2 = (|a5);
  assign y3 = (&((~(~|(~$signed($unsigned(($unsigned(a0)!==(a3)))))))!=(|$unsigned((6'd2 * (p12<a1))))));
  assign y4 = ((($signed(a3)===(b0!=b2))>>>($unsigned(p8)<<(4'd2 * b2))));
  assign y5 = (~|{{(~(b1-b2)),((~^p14)<={p9,p0})},({(b2&b5),{b1}}==={b2,b5,a1})});
  assign y6 = ((5'sd7));
  assign y7 = (a1>>a2);
  assign y8 = (+($unsigned(($unsigned((-5'sd15))/a3))==((p1>=a4)>=(b0>>a4))));
  assign y9 = (~|(-5'sd5));
  assign y10 = ((~|(&{2{p11}}))?(2'd0):(^(4'sd4)));
  assign y11 = (~|{4{p9}});
  assign y12 = ((p2&&p11)&&(~&(|p6)));
  assign y13 = (((p7+b3)>=(5'd2 * a2))?(6'd2 * (-(p6?p14:p2))):((p1?p9:a2)?(p11&&p1):(p7?p8:p16)));
  assign y14 = ((5'd22)<=((p10?a1:p14)?{a0,p15}:(p4)));
  assign y15 = (!{(p9^p17),{b2,p2,a5}});
  assign y16 = ((((p8<<<a3)>=(p6|p8))|((p15^b5)&&{b1,b0,p13}))-{(({a1,a3,b0}&&(a4|a1))===({b4}||{b2}))});
  assign y17 = (^(~&(~{(|(&$signed((~|(~|$signed(a2)))))),$unsigned(({(-(~^(p8<=p0)))}))})));
endmodule
