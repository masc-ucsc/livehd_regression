module expression_00779(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'sd15);
  localparam [4:0] p1 = ((((5'd25)>>(2'd1))<=((4'd2)^(2'sd1)))>>(4'd2 * {(5'd20),(3'd1)}));
  localparam [5:0] p2 = ((~&((2'd3)||(2'd0)))&&(-(!(2'd0))));
  localparam signed [3:0] p3 = (&(+((-3'sd0)<<{4{(5'sd15)}})));
  localparam signed [4:0] p4 = (~((4'sd2)?(4'd12):(2'sd1)));
  localparam signed [5:0] p5 = (-({3{(-4'sd4)}}===(((-3'sd3)-(4'd6))==((2'd1)!=(4'd9)))));
  localparam [3:0] p6 = (((^(-3'sd2))*((5'd31)<=(5'd4)))>=(5'd2 * ((3'd4)||(2'd3))));
  localparam [4:0] p7 = ((5'd14)?(2'd1):(4'd0));
  localparam [5:0] p8 = {4{{4{(5'd24)}}}};
  localparam signed [3:0] p9 = {{(-3'sd2),(4'd12),(-3'sd2)},{((4'd5)>>(4'sd0)),((2'd3)^(-3'sd2))},{(4'sd6),(3'd3),(2'd0)}};
  localparam signed [4:0] p10 = (({(-5'sd14),(-4'sd3)}<<<(|(2'd0)))|((|(4'sd5))!=(~(4'd0))));
  localparam signed [5:0] p11 = (-(|(((4'd5)|(4'd1))<<(3'd7))));
  localparam [3:0] p12 = {3{{3{((3'd2)>>>(3'd3))}}}};
  localparam [4:0] p13 = (((6'd2 * (2'd2))?(5'sd11):((-3'sd3)>=(3'd5)))<=(2'sd1));
  localparam [5:0] p14 = ((((5'd11)&&(-2'sd1))>={3{(-5'sd3)}})|({1{(5'sd3)}}&((-2'sd1)|(2'd0))));
  localparam signed [3:0] p15 = (-4'sd7);
  localparam signed [4:0] p16 = (5'd26);
  localparam signed [5:0] p17 = ({1{({(4'd1),(3'd0),(3'sd1)}>((-2'sd0)>=(-2'sd0)))}}>{{2{(2'd1)}},((5'sd12)|(4'd12))});

  assign y0 = {({3{b4}}?{2{p8}}:{3{a2}})};
  assign y1 = (~&(&(~|(3'd4))));
  assign y2 = (5'd2 * (~&(3'd2)));
  assign y3 = {{p9,p16,b2},(&(~&{1{p14}})),(!(-{p11}))};
  assign y4 = (4'sd3);
  assign y5 = (2'd1);
  assign y6 = $unsigned(((-(p16<a1))/a2));
  assign y7 = (5'd22);
  assign y8 = (~|((3'd0)==={{3{b4}},(4'd10)}));
  assign y9 = $signed((((p15)^(~|b4))==(3'sd1)));
  assign y10 = {3{(-3'sd1)}};
  assign y11 = (~^{b4,a1,a4});
  assign y12 = (((6'd2 * (a1?b2:a0)))-(~((b2?b3:b3)<=(+a2))));
  assign y13 = {1{((~|{4{a3}})>>>(4'd2 * (+{1{p8}})))}};
  assign y14 = ((p14?p4:p3)?(p2?p9:p6):$signed((-p14)));
  assign y15 = (2'd2);
  assign y16 = ((-p4)?{4{p6}}:{4{a3}});
  assign y17 = {({a0,a3}>={b1}),(3'd2),{(5'd12),{a4,p12},{a1,b1}}};
endmodule
