module expression_00251(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(~((-2'sd0)!=(2'sd0)))}};
  localparam [4:0] p1 = (-4'sd2);
  localparam [5:0] p2 = (((4'd4)<(-5'sd9))&&((5'sd4)>(5'sd11)));
  localparam signed [3:0] p3 = (+(((4'sd5)?(2'd3):(-4'sd5))?{(3'sd1)}:(!(3'd2))));
  localparam signed [4:0] p4 = (-5'sd6);
  localparam signed [5:0] p5 = {(((4'sd4)>(4'd9))<(&{(4'd12),(2'sd0)})),((2'd1)>{3{(2'd2)}})};
  localparam [3:0] p6 = {4{(-4'sd5)}};
  localparam [4:0] p7 = (((5'sd11)+(-2'sd1))?{4{(5'sd11)}}:((4'd13)||(3'd7)));
  localparam [5:0] p8 = ((((-3'sd1)>(5'sd9))*((2'd2)?(3'sd0):(2'sd1)))|(((5'd9)^~(5'd30))-((4'sd7)&(3'sd3))));
  localparam signed [3:0] p9 = {(-(-5'sd12)),((4'd12)?(2'sd1):(2'd3))};
  localparam signed [4:0] p10 = {{(2'd0),(4'd12),(2'd2)},((3'sd3)>>>(-5'sd2))};
  localparam signed [5:0] p11 = {3{(4'sd2)}};
  localparam [3:0] p12 = ((~&(5'd19))<<((4'd15)&(5'd24)));
  localparam [4:0] p13 = (|{1{{3{{1{(2'd0)}}}}}});
  localparam [5:0] p14 = ((3'd4)?(2'd2):(2'sd0));
  localparam signed [3:0] p15 = (-(((4'd0)?(3'sd3):(2'sd0))?{1{(4'd1)}}:{1{(2'sd1)}}));
  localparam signed [4:0] p16 = {3{(4'd2)}};
  localparam signed [5:0] p17 = ((|((5'd26)!==(5'd29)))-(|((4'sd6)&(2'sd0))));

  assign y0 = (b1&b1);
  assign y1 = (3'd7);
  assign y2 = (($signed(p16)+(3'd2))>=(-5'sd1));
  assign y3 = (2'd3);
  assign y4 = (~|($signed(({2{(a5!==a0)}}==(^(b5>a0))))^{1{{1{{2{((b5)^~(a5>a4))}}}}}}));
  assign y5 = (~((2'sd0)<<<((b0>a4)>=(&p12))));
  assign y6 = (!(~^(+{b1,b0,b0})));
  assign y7 = (!{4{(~|(|(a4+p5)))}});
  assign y8 = {2{(p12>a0)}};
  assign y9 = (-2'sd1);
  assign y10 = (4'd2 * (a1*b0));
  assign y11 = ({(&(2'd3))}<<(&(p10^p16)));
  assign y12 = (-(2'sd1));
  assign y13 = (~^b5);
  assign y14 = (b5>>>p8);
  assign y15 = ({{{b4,a5}},(b2?p0:a4),(b4<<b5)}>>(4'sd1));
  assign y16 = (-3'sd0);
  assign y17 = (((b4?a2:b1)|(p12<<p7))>((p12-a0)?(b5^~b2):{3{a5}}));
endmodule
