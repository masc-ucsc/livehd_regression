module expression_00185(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({4{(-5'sd14)}}|{2{(4'sd2)}})^(((4'd5)==(4'sd2))+(|(4'd8))));
  localparam [4:0] p1 = ((4'd10)&((4'd14)>>(((4'd8)>>(3'sd0))||{(3'sd2),(2'sd1),(3'd7)})));
  localparam [5:0] p2 = ({3{((5'sd4)==(5'sd5))}}>({4{(5'd29)}}!==(~^(~^(5'd14)))));
  localparam signed [3:0] p3 = (~^(((-4'sd5)==(5'd31))-((4'sd6)<<(2'd3))));
  localparam signed [4:0] p4 = ((~&{1{(((-2'sd1)&(5'sd0))>>(~^(5'sd7)))}})!=={2{(|(6'd2 * (3'd3)))}});
  localparam signed [5:0] p5 = ((((-(-5'sd4))%(-4'sd3))!=(4'd2))>((5'd27)*((-3'sd0)!==(-3'sd2))));
  localparam [3:0] p6 = {{(&(3'd3))}};
  localparam [4:0] p7 = {(((3'd7)?(4'sd1):(2'd2))?((-2'sd1)?(-4'sd7):(5'd30)):{(-4'sd6)}),(((4'sd2)?(5'd28):(5'd5))?((-5'sd8)>>>(3'd7)):((3'sd2)?(-3'sd3):(5'sd14))),({(3'sd1),(3'sd1),(3'd0)}+((3'd6)+(2'd0)))};
  localparam [5:0] p8 = (((5'sd3)!==(5'd29))+(5'd2 * (5'd11)));
  localparam signed [3:0] p9 = (((4'sd3)===(5'd15))%(5'd15));
  localparam signed [4:0] p10 = {2{{4{(6'd2 * (2'd0))}}}};
  localparam signed [5:0] p11 = (((5'sd2)>=(3'd6))/(3'sd1));
  localparam [3:0] p12 = (~&(((-2'sd1)>=(-2'sd1))/(-2'sd1)));
  localparam [4:0] p13 = (~^(+((!(-((2'd0)<<<(-5'sd4))))&&(((-4'sd5)&&(4'sd7))&(~(-5'sd1))))));
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = (2'd0);
  localparam signed [4:0] p16 = {1{(~^(~^(-(2'd0))))}};
  localparam signed [5:0] p17 = (((4'd2)<<<(-4'sd0))-((2'd2)===(2'd2)));

  assign y0 = ((a5+b4)!=={a2});
  assign y1 = (~|{2{{(&{b5,a2})}}});
  assign y2 = (({((p0!=p4)!=(p15-p6))}&((p4<=p9)&&{p16,p5,p11}))&&{$unsigned((6'd2 * (p12^p12))),((p5|p5)<(p16>=p15))});
  assign y3 = (3'sd2);
  assign y4 = (~|{((+(a5!==b4))!==((4'd2 * b2)-{b4,b5})),{{4{a2}},{1{(b2>>>b3)}},(~(b1-a0))}});
  assign y5 = (p15<p1);
  assign y6 = {3{$signed($signed(((-3'sd0)?(a4?b2:b4):$signed(b0))))}};
  assign y7 = (~(^({1{(2'd2)}}<<({4{p15}}<<{1{(-(a0&&a1))}}))));
  assign y8 = (~|{2{{2{((a5<=b5)&&(+a1))}}}});
  assign y9 = (((p7>p4)?((p11-p0)):(p17||p14))>(^((p4?p12:p11)?(~|(p6?p6:p6)):(p2<=p3))));
  assign y10 = (5'sd11);
  assign y11 = ((&({3{p6}}>(|p0)))<$unsigned((~(p4>>p0))));
  assign y12 = {{3{b5}},{3{b4}},{4{a4}}};
  assign y13 = (|(2'sd0));
  assign y14 = $signed({((a5&&a2)!==(5'd13)),{3{p12}},{(p13&p1)}});
  assign y15 = (!a5);
  assign y16 = (((a0?b4:p16)<{2{p6}})?{((p17>=p0)?(4'd2 * b1):{1{b4}})}:((a3>>>b3)?(a5<<<a1):(b5===b1)));
  assign y17 = $unsigned({{b2,b1,p1},{p8}});
endmodule
