module expression_00851(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(-4'sd5),(-2'sd1),(-3'sd0)};
  localparam [4:0] p1 = ((4'd0)?((4'd15)!=(3'd5)):(5'sd0));
  localparam [5:0] p2 = (({2{(5'sd4)}}?{1{(3'd1)}}:{3{(5'd7)}})?{2{((-2'sd1)?(-2'sd1):(4'd14))}}:{{(-4'sd4)},{(-5'sd3),(-2'sd1),(2'sd0)}});
  localparam signed [3:0] p3 = (5'sd12);
  localparam signed [4:0] p4 = ((&((-2'sd1)+(5'd17)))>={{(-2'sd0),(5'd26),(4'd5)},((5'd10)>>>(4'sd1))});
  localparam signed [5:0] p5 = (4'd14);
  localparam [3:0] p6 = {2{(-4'sd1)}};
  localparam [4:0] p7 = (({(2'd3),(2'd2),(4'd14)}?((-2'sd1)!=(5'd9)):(4'sd2))<{(3'd3),((4'd12)>>(2'd1))});
  localparam [5:0] p8 = (|(-{3{((-5'sd8)?(3'd1):(-5'sd13))}}));
  localparam signed [3:0] p9 = (~^(&((~|(-5'sd5))>(2'd0))));
  localparam signed [4:0] p10 = (+(4'd15));
  localparam signed [5:0] p11 = (((4'd8)?(3'd7):(2'd2))||((-2'sd1)?(5'd8):(-2'sd0)));
  localparam [3:0] p12 = (~|{4{((3'sd0)?(-5'sd3):(3'd1))}});
  localparam [4:0] p13 = ((2'sd1)==(5'd12));
  localparam [5:0] p14 = {({(2'd0),(5'd19)}==((3'sd3)?(5'd24):(4'd12))),({(2'd2),(4'sd6),(2'sd0)}?(6'd2 * (4'd15)):((-5'sd12)!=(5'd13))),(((4'd0)?(4'd11):(5'd2))?(6'd2 * (5'd2)):((5'd3)||(2'sd0)))};
  localparam signed [3:0] p15 = ((((4'sd4)?(2'sd0):(5'sd11))===(|(&(5'd30))))===(((-5'sd8)+(-3'sd2))?((-5'sd8)<=(3'sd3)):{3{(-2'sd0)}}));
  localparam signed [4:0] p16 = {2{((4'sd4)?(4'd13):(3'sd0))}};
  localparam signed [5:0] p17 = ((5'sd13)===(-5'sd12));

  assign y0 = (((!(p15?p17:p13))?$signed((~&p14)):(!$signed(a3)))<<<(~|($unsigned((^(p1?p15:b4)))&&(|(p6==p11)))));
  assign y1 = $signed((((+((b1==b5)!=(b1<<b1))))));
  assign y2 = (p4>>>b0);
  assign y3 = $unsigned(($unsigned(p16)/p7));
  assign y4 = ((2'd1)?(4'sd4):(^(-2'sd1)));
  assign y5 = $signed($signed($unsigned((|(~^((-(p9?a1:p15))<=(&(p3?p4:p11))))))));
  assign y6 = ((~^(!(&(!((b3===b2)<(&(~p4)))))))|(!(-(-((b0||a5)<<<(p0<<p1))))));
  assign y7 = {(&(&{2{a0}})),({a2,a1}===(^a2)),{4{a1}}};
  assign y8 = (-3'sd3);
  assign y9 = (a1?p1:p14);
  assign y10 = ((~&{(b5||p17)})||(~&(b5^~p17)));
  assign y11 = (!((|p10)||(^p8)));
  assign y12 = (({(b5?p8:p0),{b4,b2}})<(~^({3{p17}})));
  assign y13 = (b1?b2:p7);
  assign y14 = (&(~(~^(-5'sd6))));
  assign y15 = (-(|((-(~|(2'd3)))<((-5'sd8)?{3{b5}}:(!(&b0))))));
  assign y16 = (((a5?p0:b1)+($signed(a2)!==(a1!=b3)))>$unsigned(((!(~|p11))+(2'd0))));
  assign y17 = (&a3);
endmodule
