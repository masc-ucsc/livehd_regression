module expression_00371(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(((2'd2)&&(4'd3))&((4'd0)+(-4'sd0)))}};
  localparam [4:0] p1 = {(((2'sd1)===(4'd0))<<<{(3'd1)}),({(3'd1),(-3'sd3),(5'sd3)}=={(-4'sd3),(-3'sd0)})};
  localparam [5:0] p2 = (!((3'd5)?(-2'sd1):(-5'sd3)));
  localparam signed [3:0] p3 = ({((2'd1)>>>(5'd5)),(+(-4'sd7)),(5'sd7)}==(((3'd7)&&(2'd2))-((3'd0)>=(5'd14))));
  localparam signed [4:0] p4 = {(5'd3)};
  localparam signed [5:0] p5 = (5'sd3);
  localparam [3:0] p6 = (({(-3'sd3)}-{(2'sd1),(3'd5)})<<<(((2'd2)<<(-3'sd1))|((5'd7)&&(3'sd0))));
  localparam [4:0] p7 = ((((-3'sd2)^(2'd3))!=((-5'sd6)==(4'sd7)))<(((3'sd1)%(-5'sd6))-((2'd1)|(5'd2))));
  localparam [5:0] p8 = (&(~&(-2'sd1)));
  localparam signed [3:0] p9 = {((5'd8)^(((2'd1)>(4'd9))!=={(2'd0),(5'd4)}))};
  localparam signed [4:0] p10 = ({(3'd1),{(5'sd15),(4'd12),(-3'sd0)},(+(2'd0))}<<<(-3'sd1));
  localparam signed [5:0] p11 = {{4{(-2'sd0)}},{(3'sd2),(2'd3)}};
  localparam [3:0] p12 = {({{(-4'sd0),(5'd27),(2'd3)},((4'sd6)||(2'd1))}!==(((4'd9)>(4'sd3))&((5'd1)|(5'd12))))};
  localparam [4:0] p13 = (-(5'd2 * ((5'd21)!==(3'd3))));
  localparam [5:0] p14 = (3'sd2);
  localparam signed [3:0] p15 = ({((5'd18)==(5'd25)),((3'sd0)==(3'd0)),(4'd2)}^{{(-4'sd5),(4'd2)},(-2'sd1),((-4'sd3)||(3'd3))});
  localparam signed [4:0] p16 = (-{(-3'sd3),(5'sd11)});
  localparam signed [5:0] p17 = {(2'sd1),(+(!(~&((4'sd0)!=(3'd4)))))};

  assign y0 = (4'd1);
  assign y1 = (~&(((+(~^(p2^~a4)))>((b3<p7)||(b1||a2)))^(^(~|((+(a3===b3))==(p16+p11))))));
  assign y2 = ((a2!=a0)?(~(b1&a3)):($unsigned(b4)));
  assign y3 = ({3{{1{a1}}}}>{4{(-2'sd0)}});
  assign y4 = $unsigned(({2{((b0===a2)<{3{b0}})}}!=($unsigned((5'd2 * p12))<<<{3{p2}})));
  assign y5 = (~p13);
  assign y6 = (b1===a0);
  assign y7 = ((p16|p7)?{(p10?p17:a5)}:(b2^~p8));
  assign y8 = (-5'sd0);
  assign y9 = (((~|p13)?{2{p11}}:(p3-p5))&&(+({3{p4}}?(p6>>p6):{3{b1}})));
  assign y10 = {(p17|p5),(p9^p10),(p8==p3)};
  assign y11 = (|((~^$signed((~|a5)))&((^p8)/b3)));
  assign y12 = ({2{a4}}?(a5&b4):(a4?b2:b1));
  assign y13 = {2{(6'd2 * p12)}};
  assign y14 = ({$unsigned(b1),$unsigned(p10)});
  assign y15 = (^(p3?p7:p11));
  assign y16 = (((^(5'd2 * (b1?a1:a0))))<<<((a3)?(+a1):$unsigned(a5)));
  assign y17 = (-{{{b1,b0,a0},{p5,a3}},({p14,b1}<=(b2?b3:a3))});
endmodule
