module expression_00184(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(2'sd1)};
  localparam [4:0] p1 = {(!{3{(3'd1)}}),{3{(3'd2)}}};
  localparam [5:0] p2 = {(((5'd24)==(3'sd0))?{(-2'sd0),(-4'sd4)}:((3'd6)||(5'd8)))};
  localparam signed [3:0] p3 = ((2'd1)?(-3'sd1):(-2'sd0));
  localparam signed [4:0] p4 = (4'd2);
  localparam signed [5:0] p5 = (((2'd1)?(3'd0):(-3'sd1))?((5'sd11)?(3'sd1):(-2'sd0)):((3'sd3)>>>(3'd0)));
  localparam [3:0] p6 = (~|({(|{((2'd3)>=(-4'sd2))})}-(~|{(2'd0),(-2'sd0),(3'd5)})));
  localparam [4:0] p7 = (2'sd1);
  localparam [5:0] p8 = ((3'd7)-(-3'sd3));
  localparam signed [3:0] p9 = {4{(5'd17)}};
  localparam signed [4:0] p10 = ({((2'd3)+(-3'sd3))}>=(4'd11));
  localparam signed [5:0] p11 = {((((2'sd0)?(3'd7):(5'd1))?(4'd2 * (2'd1)):((5'sd9)?(3'd6):(-2'sd0)))||(((3'd3)?(5'd24):(-2'sd1))?((-3'sd3)>>(-5'sd6)):{(-5'sd10),(3'sd0)}))};
  localparam [3:0] p12 = (5'd24);
  localparam [4:0] p13 = (2'd3);
  localparam [5:0] p14 = ((((5'd24)|(5'd17))!==((4'd11)?(4'sd2):(-2'sd0)))-(((4'sd1)+(5'sd4))<<<((2'd1)<<(-5'sd10))));
  localparam signed [3:0] p15 = ((((5'sd2)|(-2'sd1))?((3'sd1)?(5'd13):(4'sd7)):{(2'd0)})^~(((-5'sd8)>>>(2'sd1))&{(2'd2),(2'sd0),(-5'sd9)}));
  localparam signed [4:0] p16 = (-2'sd0);
  localparam signed [5:0] p17 = (~|(+(2'd3)));

  assign y0 = (2'd1);
  assign y1 = (&(!(-((~b4)&(~^p11)))));
  assign y2 = {(-$unsigned((b5))),{(~|(b0?a0:p16))},{{(a1===b1)}}};
  assign y3 = (~^p6);
  assign y4 = (4'd9);
  assign y5 = {1{({2{{$unsigned({a0,b5,b4}),{a4,a1}}}})}};
  assign y6 = {{(a2!==b3),(b4!==a0),(p11)},({4{p10}}!=(~a4)),$unsigned(((p17||b2)>=$signed(p8)))};
  assign y7 = ((((a1||p9)^(p6<<<p8))|(2'd2))=={3{(a4&&b3)}});
  assign y8 = ((~|p16)?(p10?p17:p6):(&p14));
  assign y9 = {4{(p10>p2)}};
  assign y10 = (~^({a3}<<<{p5,a4}));
  assign y11 = (3'd7);
  assign y12 = (-({1{(({1{a2}}||(a1<<<b5))<<<((-b2)>={1{b4}}))}}<<<{2{((a5!==b1)<<(b5+b1))}}));
  assign y13 = ((p0?p16:b4)?(-2'sd1):(-3'sd1));
  assign y14 = (|{4{(|(b3<<<a3))}});
  assign y15 = ((+{{a5,b2},(b5^a1),(b3!=b0)})>>>({{(a2>=a1)}}===((5'd26)^(a5!=a1))));
  assign y16 = ($unsigned((b3-a3))!==(-4'sd2));
  assign y17 = ((b3==b2)?(b2>>b3):(b5!=a3));
endmodule
