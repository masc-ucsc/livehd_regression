module expression_00388(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (|((~|(&{(5'd22)}))|{4{(3'd6)}}));
  localparam [4:0] p1 = ({((5'd12)&&(2'd3))}===((3'd1)|(4'sd5)));
  localparam [5:0] p2 = (5'd28);
  localparam signed [3:0] p3 = ((((-3'sd3)|(4'sd7))+((-3'sd2)^(5'd12)))<=(-5'sd5));
  localparam signed [4:0] p4 = (^{4{(3'd3)}});
  localparam signed [5:0] p5 = {1{{2{(2'sd0)}}}};
  localparam [3:0] p6 = {{1{({3{{3{(2'sd0)}}}}^~{({(4'd8)}&{4{(5'sd15)}})})}}};
  localparam [4:0] p7 = (-2'sd1);
  localparam [5:0] p8 = ((|{3{(5'sd9)}})<<<(4'd2 * (5'd6)));
  localparam signed [3:0] p9 = {4{(2'd1)}};
  localparam signed [4:0] p10 = (((3'sd1)&(3'sd1))?{1{(4'd1)}}:{3{(-3'sd3)}});
  localparam signed [5:0] p11 = (^(-({2{{1{(3'd2)}}}}+(~(~|((3'd2)<(3'd6)))))));
  localparam [3:0] p12 = {1{{1{{((3'd6)?(-3'sd0):(4'sd5))}}}}};
  localparam [4:0] p13 = (4'd3);
  localparam [5:0] p14 = (-(^{{(2'd1),(5'sd5),(5'sd12)}}));
  localparam signed [3:0] p15 = ((3'sd0)<<(|{(3'sd0),(3'd3),(-5'sd14)}));
  localparam signed [4:0] p16 = ((2'sd1)||(-3'sd0));
  localparam signed [5:0] p17 = (~&{(6'd2 * (5'd2 * (3'd7))),{4{(3'sd1)}}});

  assign y0 = (p13^~b4);
  assign y1 = ({({4{a1}}<<<{3{b1}}),((a1<=a3)+(a0&&a0))}<=(((a3+b3))&&({4{a4}})));
  assign y2 = (~|((|p10)>>(p10<<<p7)));
  assign y3 = ({(p12-p3),{3{p16}},(-{4{p0}})}>>{{((|p12)-$signed(p15)),{2{(p4&&p11)}}}});
  assign y4 = ((~|(~{p16,b2}))<={4{a0}});
  assign y5 = {4{$signed(a0)}};
  assign y6 = (5'd27);
  assign y7 = (^(~&(((b2>>b0)>(a1?b5:b4))<<<((a0&a3)-(p10>=p5)))));
  assign y8 = ((-5'sd12)>(3'sd3));
  assign y9 = (4'd2 * (~^(p12-b1)));
  assign y10 = ((p13^~p9)?{{p9,b3,p3}}:$unsigned((p10>=p2)));
  assign y11 = {2{{{(a4)},{a3,b3,a2},(p1<=a2)}}};
  assign y12 = (4'd15);
  assign y13 = ((~(&{4{p8}}))?(|(~&(p10?a5:b0))):{4{(~b3)}});
  assign y14 = (~|((4'sd2)>>((p17<p0)<<(p17*p0))));
  assign y15 = (^({3{p0}}||(-5'sd7)));
  assign y16 = {{{3{$unsigned($signed((b3)))}}}};
  assign y17 = {1{{4{{3{{p8}}}}}}};
endmodule
