module expression_00194(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(^{{3{(2'd0)}},((5'sd5)?(4'd15):(-5'sd10)),((5'd10)?(-3'sd1):(-5'sd15))}));
  localparam [4:0] p1 = ((((2'sd0)&(2'sd1))&&((2'd3)^~(4'sd6)))?{4{(3'd2)}}:{4{(-4'sd4)}});
  localparam [5:0] p2 = (-((~^((!((-2'sd0)<<(3'sd3)))<(~((-5'sd12)||(-5'sd15)))))<(~&((!(-(4'sd3)))<<((-3'sd0)&&(-3'sd3))))));
  localparam signed [3:0] p3 = (-4'sd0);
  localparam signed [4:0] p4 = (5'd30);
  localparam signed [5:0] p5 = (((5'sd12)?(5'sd9):(-4'sd5))>>((-2'sd1)<<<(-5'sd2)));
  localparam [3:0] p6 = {1{{2{((-2'sd0)?(5'sd9):(3'd6))}}}};
  localparam [4:0] p7 = ((!(5'd0))?((-2'sd0)>(-2'sd1)):(-2'sd0));
  localparam [5:0] p8 = (((3'sd2)/(5'd22))?((-5'sd7)?(3'sd1):(-3'sd2)):((-5'sd1)>=(2'sd0)));
  localparam signed [3:0] p9 = (~&({(-{(2'd1),(2'sd0),(2'd3)})}>=((&((2'sd1)&(5'sd6)))-(-4'sd7))));
  localparam signed [4:0] p10 = (|(~^(((3'd2)|(5'sd12))>>(-(5'sd4)))));
  localparam signed [5:0] p11 = ((-5'sd13)||(4'd10));
  localparam [3:0] p12 = ({((4'd9)>=(-4'sd2)),{(4'd10),(-4'sd1)},((4'sd1)||(-3'sd1))}>>>{(4'd14),(-(2'sd0)),((-5'sd6)&(5'sd15))});
  localparam [4:0] p13 = ({((5'd13)?(4'sd5):(-4'sd2))}?((+(5'd2))?((-3'sd3)?(3'd7):(-3'sd2)):((2'd0)<(-3'sd2))):(-({(-3'sd1)}>>>((3'sd1)>>>(5'd21)))));
  localparam [5:0] p14 = (-((^(2'd3))||((~^(-2'sd1))^(-(5'd9)))));
  localparam signed [3:0] p15 = (~((((-3'sd1)<=(4'd15))>(^(3'sd0)))?(((-2'sd0)<(2'sd1))+((3'sd2)^(4'd12))):({(5'd13)}?((5'sd4)>>>(-3'sd0)):((5'd29)?(5'd9):(4'sd4)))));
  localparam signed [4:0] p16 = {3{{1{(4'd7)}}}};
  localparam signed [5:0] p17 = (~{1{(5'd14)}});

  assign y0 = (((b5==b3)<={1{b4}})?((b1>>>p4)?{4{b1}}:(-p17)):{3{(p1+b2)}});
  assign y1 = (3'sd0);
  assign y2 = (p17<<b0);
  assign y3 = $signed(((((-3'sd3))>(2'sd0))+((p12-p7)-$unsigned((p15?p14:p4)))));
  assign y4 = (&(~({3{(-p12)}}|{2{(!{4{p5}})}})));
  assign y5 = {({p10,p1,a2}&(p13&p9))};
  assign y6 = ((-3'sd2));
  assign y7 = (6'd2 * b0);
  assign y8 = ((5'sd4)?$unsigned((6'd2 * {2{a0}})):((4'd2)?(a3<<a3):$signed(b5)));
  assign y9 = (({p8,p17,p9}-(p11&&p2))^~({p0,p3,p7}^~(|(p9==p16))));
  assign y10 = (4'sd4);
  assign y11 = ((b5||a0)?(a5!==a2):(|a4));
  assign y12 = $signed({1{{4{(+(-(~&p3)))}}}});
  assign y13 = $unsigned(((&(2'sd0))));
  assign y14 = ((p8^~p15)?{p8,a5}:{1{p17}});
  assign y15 = $unsigned((~|{1{{{p12,p10},{b1}}}}));
  assign y16 = ({{{2{{$signed(a3),(b1)}}},{4{(a2)}}}});
  assign y17 = {4{(~&p10)}};
endmodule
