module expression_00700(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'sd1);
  localparam [4:0] p1 = (-2'sd0);
  localparam [5:0] p2 = (((5'd25)?(2'd3):(3'd1))?(4'sd2):((4'sd1)?(3'd1):(5'sd7)));
  localparam signed [3:0] p3 = ({{1{((3'd5)<=(4'd3))}}}>>>{4{(4'd10)}});
  localparam signed [4:0] p4 = (-(-2'sd0));
  localparam signed [5:0] p5 = ({1{{4{(3'sd2)}}}}>=((-4'sd1)?(5'sd1):(4'd4)));
  localparam [3:0] p6 = ({(&{2{(2'sd1)}}),(^{2{(2'sd1)}}),(|((3'd7)==(4'sd1)))}|{{4{(4'sd5)}},(|((5'd10)!=(5'sd5)))});
  localparam [4:0] p7 = (~(!(-2'sd0)));
  localparam [5:0] p8 = (((4'sd6)^~(5'sd13))*((3'd5)<=(3'sd1)));
  localparam signed [3:0] p9 = ((-(~^(~(~&(2'd1)))))<<(+{1{(~{3{(5'd17)}})}}));
  localparam signed [4:0] p10 = (~^((~((4'sd6)?(-4'sd6):(3'sd1)))?(3'd5):({(-4'sd1),(5'd31),(4'd15)}?{(5'd3),(-5'sd14)}:(-3'sd3))));
  localparam signed [5:0] p11 = (((4'd1)?(4'd9):(3'd0))>={(4'sd2),(4'd3),(2'd2)});
  localparam [3:0] p12 = (-(^(-2'sd1)));
  localparam [4:0] p13 = (~^{(&(-3'sd3)),(~^(2'd1)),(~^(3'sd1))});
  localparam [5:0] p14 = (6'd2 * {4{(5'd31)}});
  localparam signed [3:0] p15 = (+((~(3'sd3))<<((2'sd1)!=(3'sd2))));
  localparam signed [4:0] p16 = (~^(|(((3'sd3)-(5'd18))|(|(2'd2)))));
  localparam signed [5:0] p17 = ({3{(&(5'd3))}}>>(((-5'sd4)?(5'd22):(3'd5))^((4'sd6)?(4'd5):(5'sd13))));

  assign y0 = (((b5+b2)-{a1,a0})-((a1^p0)^~$signed($signed(a1))));
  assign y1 = (!(((a0^b0)!==(~&(a0?b5:a2)))<<(5'd2 * (p7?p7:p12))));
  assign y2 = ((~&((a1<p5)^~(5'sd10)))>=((b2&&b0)||(~p17)));
  assign y3 = ({2{{4{p6}}}}<<{{1{b3}},{a0},$unsigned(p15)});
  assign y4 = (+({3{(~&b2)}}&&{2{(b0-b3)}}));
  assign y5 = (-(~^(p3?a3:a2)));
  assign y6 = (2'd2);
  assign y7 = (~|({4{a4}}!==(~(b1==a2))));
  assign y8 = (5'sd3);
  assign y9 = ((~(b5*a0))>>>((a4^~p9)==(a1?p9:b2)));
  assign y10 = (~^(~^({2{(&a4)}}?((b3+b1)>>(~b3)):(-5'sd9))));
  assign y11 = ((a5!=p1)*(p13^~a2));
  assign y12 = $signed((-4'sd1));
  assign y13 = ((!(((2'd0)!==(a5?a0:a3))!==({3{a5}}^(~&b3))))>=(((b0?p2:b5)<(a0+p6))-({b5,a4}|{b1,p12,a0})));
  assign y14 = (6'd2 * (b0>>p1));
  assign y15 = ({{a2,a1},(p17<<<a0),(p3||b2)}<<<((p4?b3:a1)?(a0-b2):{b0,p3}));
  assign y16 = (p9?p5:p4);
  assign y17 = (+$signed((~&(|{2{(-{((~^{p17}))})}}))));
endmodule
