module expression_00383(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(((5'd3)>(-2'sd0))+((-3'sd0)!=(3'd5)))}};
  localparam [4:0] p1 = (~(~&(&(~&(+(~(~^(~(|(2'sd0))))))))));
  localparam [5:0] p2 = (|{1{(4'sd4)}});
  localparam signed [3:0] p3 = (-3'sd3);
  localparam signed [4:0] p4 = (((2'sd0)>>>((4'sd1)^~(4'd14)))?((3'sd1)!=((4'sd7)?(2'd3):(3'd2))):(((5'd24)>>>(4'd4))^((4'sd6)%(4'sd2))));
  localparam signed [5:0] p5 = (4'd6);
  localparam [3:0] p6 = (3'd0);
  localparam [4:0] p7 = ((~^(^(~|(^{(~{4{(2'd2)}})}))))<<<(&(|(((4'd15)<=(4'd8))+(&{3{(5'sd10)}})))));
  localparam [5:0] p8 = (({(-2'sd1)}|((3'sd3)||(5'd22)))&({(2'd3)}!=(3'd7)));
  localparam signed [3:0] p9 = (-2'sd1);
  localparam signed [4:0] p10 = {2{{2{{1{(4'd2 * (4'd6))}}}}}};
  localparam signed [5:0] p11 = ({1{{((3'd5)!==(-2'sd1)),(4'd2 * (5'd3))}}}>=(({2{(2'd3)}}!==((-2'sd0)|(2'sd1)))^{{3{(5'd6)}}}));
  localparam [3:0] p12 = {4{{1{{2{(4'd3)}}}}}};
  localparam [4:0] p13 = (-3'sd3);
  localparam [5:0] p14 = ((({(4'sd1)}>{(3'sd0),(5'd14)})=={(5'd7),(4'sd7),(3'd0)})<<(4'd2 * ((3'd5)|(5'd14))));
  localparam signed [3:0] p15 = ((({(4'd5),(4'd7)}<<<((-4'sd4)!=(2'd0)))>=(((5'd19)+(2'd2))>((5'sd7)||(5'sd10))))===(((-(4'd4))|(^(2'sd0)))-(!((5'd11)<<(4'd10)))));
  localparam signed [4:0] p16 = (3'd7);
  localparam signed [5:0] p17 = ((2'sd1)!==(5'd19));

  assign y0 = ((((p3+p4)!={1{p17}})>>((p2<p0)>=(p13>=p8)))>>{3{(p14?b3:p7)}});
  assign y1 = ({2{(p8&&p4)}}>>>((p0<<p0)==(4'd2 * p13)));
  assign y2 = ((b0?b4:p5)?(|b5):(5'd0));
  assign y3 = $unsigned(((-((+(-p7))))?{2{{2{p7}}}}:(-4'sd3)));
  assign y4 = ((|(~^$signed($signed(p10)))));
  assign y5 = {{{b5,b4,a1}}};
  assign y6 = (5'd17);
  assign y7 = (2'sd1);
  assign y8 = ((&(5'd2 * a1))&&(b2<<b1));
  assign y9 = (5'd0);
  assign y10 = (|(^((6'd2 * p13)<(3'sd1))));
  assign y11 = (~{2{((a4?p7:p7)?(p16?a4:a1):(b5?a3:p7))}});
  assign y12 = $unsigned((a5?b1:a0));
  assign y13 = (((a0==a0)!=(a2<<b0))>=((b5|b3)>=(b4===b0)));
  assign y14 = $signed((~^$unsigned({{p7},$signed(p16),(|b3)})));
  assign y15 = (~|$signed($signed((({4{p14}}<=$unsigned((~^(p17>>>a4))))=={1{(^((4'd2 * {2{p0}})))}}))));
  assign y16 = (^(((~(~&a0))/p0)|((p7==a1)|(a4>b3))));
  assign y17 = ({({p17,p7,p7}+(p12!=p10))}||{((p17<p14)>>>{p6,p0,p10})});
endmodule
