module expression_00260(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{{2{(-5'sd10)}}}};
  localparam [4:0] p1 = {1{(-3'sd0)}};
  localparam [5:0] p2 = (2'd0);
  localparam signed [3:0] p3 = (-(~^(3'sd2)));
  localparam signed [4:0] p4 = (~((4'd2 * {(3'd4),(4'd7),(4'd2)})+(-3'sd1)));
  localparam signed [5:0] p5 = {4{(|{3{(-4'sd3)}})}};
  localparam [3:0] p6 = {1{{1{(&{2{(~&(-3'sd0))}})}}}};
  localparam [4:0] p7 = (+(-({2{(5'd31)}}?((-4'sd2)-(5'd1)):((4'sd7)<=(4'sd2)))));
  localparam [5:0] p8 = (((-5'sd3)&(4'sd5))>=(4'd2 * (4'd8)));
  localparam signed [3:0] p9 = ((|(~|(&(-3'sd2))))===(((3'd3)>(5'd9))<((4'd7)==(4'sd6))));
  localparam signed [4:0] p10 = (((4'sd1)<(5'd21))?((-5'sd3)^~(-4'sd0)):((5'd1)+(3'd3)));
  localparam signed [5:0] p11 = (|{3{{2{{4{(2'd2)}}}}}});
  localparam [3:0] p12 = (&((-2'sd1)*(-2'sd0)));
  localparam [4:0] p13 = (({4{(3'd5)}}?((2'd2)||(2'd3)):((4'd9)||(2'sd0)))!=(((-4'sd3)+(5'sd5))?(-4'sd2):{4{(-3'sd1)}}));
  localparam [5:0] p14 = (((5'd4)<=(2'd3))&{(5'sd14),(3'd5),(5'sd3)});
  localparam signed [3:0] p15 = ((~^(~|(-5'sd2)))>>(^(!(4'd6))));
  localparam signed [4:0] p16 = (((2'sd1)%(4'd7))?((4'd14)>>(4'd15)):((3'd5)===(2'sd0)));
  localparam signed [5:0] p17 = (~{2{{1{{4{(4'd10)}}}}}});

  assign y0 = (4'd2 * (p6?p8:p8));
  assign y1 = {2{(^((a5?p0:a4)?(b1&b1):(~^p2)))}};
  assign y2 = ((-(^$signed(((a0^b4)<<(3'd0)))))!=$unsigned(($unsigned(a4)?(a4%a0):(!b4))));
  assign y3 = ((|(&(~|$unsigned(($signed({$unsigned(p5)})))))));
  assign y4 = {3{(~&(3'd5))}};
  assign y5 = (^((+(!{(&b5)}))>((b4>a5)&&(4'sd0))));
  assign y6 = ((p6|p4)?(a2||b1):(~&(b4!==a4)));
  assign y7 = (4'd1);
  assign y8 = ((2'sd1)^{(5'd26)});
  assign y9 = {4{(b0&&b2)}};
  assign y10 = (~(~$signed((!(!((-2'sd0)%p10))))));
  assign y11 = ((b4>p4)?(~p5):(p17==a0));
  assign y12 = $unsigned((((b1<b0))>>>((p15!=a1)/p3)));
  assign y13 = (~&((b3<=b0)<(a2)));
  assign y14 = (~^(~|($signed((~|{3{p3}}))?{1{((p15?p5:b2)<<(p15<<<p12))}}:{1{(p14?b5:p13)}})));
  assign y15 = ({({p3,p1}>=(a4<p2)),{(p0?p5:p3)}}!=(((p15+p3)?(p5?p11:a1):(p7<<b1))+({p6,b5,b4}==(a2<<<p11))));
  assign y16 = (~&((2'd3)>(~|(2'd3))));
  assign y17 = (2'd2);
endmodule
