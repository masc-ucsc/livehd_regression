module expression_00058(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd6);
  localparam [4:0] p1 = {1{{2{{({3{(-5'sd5)}}||(~|{(3'd0),(3'sd0),(-2'sd0)}))}}}}};
  localparam [5:0] p2 = (((-(-4'sd4))?((3'sd3)==(3'd5)):(3'd3))^~((3'sd2)?{(-3'sd3),(2'd1)}:((-5'sd14)?(4'd8):(3'd5))));
  localparam signed [3:0] p3 = (({3{(-5'sd2)}}?((3'd6)?(-4'sd0):(-2'sd0)):((4'd10)!==(3'sd2)))?{1{{2{((3'd3)^~(3'd3))}}}}:({2{(-3'sd3)}}?((3'd1)==(-4'sd6)):((4'd9)|(4'd13))));
  localparam signed [4:0] p4 = (((-5'sd13)<<<(4'sd7))!==(&(4'd12)));
  localparam signed [5:0] p5 = ((-((3'sd3)!=(2'd3)))?{2{(-4'sd1)}}:((5'sd9)?(5'sd15):(5'sd6)));
  localparam [3:0] p6 = {(2'sd0),(-3'sd2),(3'd3)};
  localparam [4:0] p7 = {2{{4{((4'sd1)?(-4'sd0):(4'sd4))}}}};
  localparam [5:0] p8 = ((2'd2)===(-3'sd1));
  localparam signed [3:0] p9 = (((2'sd1)%(4'd9))*((-4'sd2)?(4'sd3):(5'sd0)));
  localparam signed [4:0] p10 = (4'd13);
  localparam signed [5:0] p11 = ((~(4'sd0))>>>(-(2'd1)));
  localparam [3:0] p12 = (-2'sd0);
  localparam [4:0] p13 = (2'sd1);
  localparam [5:0] p14 = (4'd2);
  localparam signed [3:0] p15 = {2{{4{{(-2'sd1),(4'sd5)}}}}};
  localparam signed [4:0] p16 = {4{{4{(-3'sd1)}}}};
  localparam signed [5:0] p17 = (((5'd16)?(5'd8):(3'd5))?(!{2{(3'sd3)}}):{1{((5'sd13)&(2'd0))}});

  assign y0 = {4{((p9<<p17)-(p5>a0))}};
  assign y1 = (-3'sd0);
  assign y2 = ((p9?p1:p9)?(p4-a5):(p7-p0));
  assign y3 = ((2'd3)+((5'd15)<(2'd3)));
  assign y4 = $unsigned({4{({p7,p8}>(p1?p14:b1))}});
  assign y5 = ((^(&(~^p14)))?(p14?p3:p6):(p14?p9:p3));
  assign y6 = ({(~&(p0?a1:p14)),{(p1?a3:p17)}}?(5'd18):(-(|(^(3'sd3)))));
  assign y7 = (-(a5>>>a5));
  assign y8 = (((&a3)?(a1|p10):(+a1))&&((b0*b1)<(~(6'd2 * b2))));
  assign y9 = $unsigned($unsigned($unsigned((^b4))));
  assign y10 = ((a5-b1)>=(a1!==a0));
  assign y11 = (((b2^p13)-(p11&&p7))>>>((b5+p16)?{p13,a5,p14}:(~&p0)));
  assign y12 = ((p6+a5)||{1{(p15)}});
  assign y13 = (((6'd2 * p8)>(b3+b4))+((p9-p9)>>>(~{2{b3}})));
  assign y14 = (~|(5'd22));
  assign y15 = (p9|p17);
  assign y16 = ((3'd2)<=((4'sd4)%p13));
  assign y17 = {((b5==a1)<{b0,b0}),((~b1)||(a0>>>b0))};
endmodule
