module expression_00352(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&{{1{{3{(3'd4)}}}},{((-4'sd1)||(-5'sd8)),{4{(-2'sd0)}},{(4'd7),(3'sd3),(5'd18)}},{2{{(3'd7),(-4'sd1)}}}});
  localparam [4:0] p1 = (-3'sd0);
  localparam [5:0] p2 = ({2{(~&{1{(5'd24)}})}}||(~(^(|(&{1{(5'd14)}})))));
  localparam signed [3:0] p3 = (6'd2 * (-(!(3'd5))));
  localparam signed [4:0] p4 = {(4'd2 * ((5'd6)-(2'd2)))};
  localparam signed [5:0] p5 = ((((4'd11)>>(-4'sd3))!==((5'd3)?(-2'sd1):(3'd1)))>>>(((5'd14)>(5'd0))!==((3'd4)<(3'sd1))));
  localparam [3:0] p6 = ((^(3'sd3))>>(~^(-4'sd2)));
  localparam [4:0] p7 = ((~|(5'd20))-((5'd27)?(2'd2):(4'd10)));
  localparam [5:0] p8 = ((2'd2)?(4'd15):(4'd6));
  localparam signed [3:0] p9 = ((^(^(4'd6)))?{1{((4'sd2)?(5'd20):(2'sd1))}}:(+(~(-5'sd11))));
  localparam signed [4:0] p10 = ((~^(5'sd6))^((5'd25)>=(-4'sd2)));
  localparam signed [5:0] p11 = (4'd8);
  localparam [3:0] p12 = (2'sd0);
  localparam [4:0] p13 = {((5'd10)?(-2'sd1):(3'd2)),((3'd0)?(3'd2):(-3'sd0))};
  localparam [5:0] p14 = {{4{(3'sd2)}},{{(3'sd0),(5'd13)},((5'd28)?(5'd4):(4'd6)),{1{(4'sd6)}}}};
  localparam signed [3:0] p15 = (3'sd0);
  localparam signed [4:0] p16 = (((-2'sd1)<=(5'd21))<((3'sd0)?(4'd1):(2'd3)));
  localparam signed [5:0] p17 = (((3'd5)<<(-5'sd12))!==((5'd23)<<<(4'd4)));

  assign y0 = (-4'sd0);
  assign y1 = (2'sd1);
  assign y2 = (5'd10);
  assign y3 = (a3+b5);
  assign y4 = {2{{3{p6}}}};
  assign y5 = {4{{{b2,a4},(p1>p14)}}};
  assign y6 = (((b3?p5:p12)+(a3&b1))<{(5'sd5),(p11>>>a5)});
  assign y7 = ({{a1,b0,p5}}&&{b4,a4,a1});
  assign y8 = (~&(((b5?p6:a2)>>>(p1?p8:b5))?(^(5'd2 * (!b1))):(^(a3?a5:b2))));
  assign y9 = ({3{{3{a2}}}}?{4{a4}}:((a3?b0:b2)^(-a1)));
  assign y10 = ((4'd2 * {a0})<<((a0^p17)|(a2?b0:b1)));
  assign y11 = ({((p13<<<p16)<<<{p12,p11,p4}),((6'd2 * p7)<<<(p11|p9))}>=(((p5-p13)+{p7})>>{{(p3+p13),{p1,a5,p16}}}));
  assign y12 = {1{(({1{(b4+p17)}}<=(&(p14+b4)))&&((b1?a5:a4)>(~|{3{p6}})))}};
  assign y13 = ($signed($unsigned((+(|((b1?b1:b3)!==((b0<=b1)))))))<(($unsigned((~(p2?p0:p15)))^((4'd2 * p12)&&(p14-p15)))));
  assign y14 = (&(!((-((4'sd5)>(a5<b0)))+(|(^((|(|p15))^(p12|p0)))))));
  assign y15 = ({1{($unsigned($signed({a3}))||{1{({2{b4}})}})}}<=(($unsigned(b5)>>(a4))<=({2{p11}}<<(a2<a3))));
  assign y16 = {3{(-5'sd14)}};
  assign y17 = (3'd5);
endmodule
