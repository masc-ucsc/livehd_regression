module expression_00241(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd2);
  localparam [4:0] p1 = (((~^(-2'sd1))?((3'd4)>>(-3'sd1)):(+(2'sd0)))?(((4'd12)&(3'sd3))*((2'd2)?(3'sd1):(5'd4))):((+(4'd11))==((3'sd2)&(3'd1))));
  localparam [5:0] p2 = ((~(~|(((2'd3)^(-2'sd1))>>>(~(+(5'sd6))))))&(4'd2 * (|((2'd3)^~(5'd3)))));
  localparam signed [3:0] p3 = (~|{{3{(~(-2'sd0))}},{4{(5'sd7)}}});
  localparam signed [4:0] p4 = (((5'd26)<<(4'sd1))+(5'sd14));
  localparam signed [5:0] p5 = ((3'sd0)?({3{(-4'sd7)}}?(&(3'd2)):((-4'sd1)==(3'd7))):{2{{(2'sd0)}}});
  localparam [3:0] p6 = {(2'd2),(-3'sd0),(5'd19)};
  localparam [4:0] p7 = (-3'sd3);
  localparam [5:0] p8 = (2'sd0);
  localparam signed [3:0] p9 = (5'sd13);
  localparam signed [4:0] p10 = ((~&((4'sd1)<(-4'sd2)))%(5'sd4));
  localparam signed [5:0] p11 = (5'sd10);
  localparam [3:0] p12 = (!(-5'sd12));
  localparam [4:0] p13 = {(((5'd27)>>>(3'd1))>{1{(2'd2)}}),({(2'd2)}>>>{2{(-3'sd3)}})};
  localparam [5:0] p14 = ((((3'sd3)?(-5'sd10):(4'd2))^~((3'd7)-(5'd21)))<<<(((-3'sd0)?(-5'sd13):(5'sd15))^~((-4'sd3)?(4'd4):(4'd1))));
  localparam signed [3:0] p15 = {{((3'sd2)>(5'sd15))},((3'sd1)|(5'd24))};
  localparam signed [4:0] p16 = (~&(2'd2));
  localparam signed [5:0] p17 = {((-5'sd15)|(3'sd2)),(~^(2'sd1)),((-2'sd1)<<(5'd26))};

  assign y0 = (-5'sd0);
  assign y1 = (^(-4'sd1));
  assign y2 = {4{({3{p5}}>>(p11==p10))}};
  assign y3 = $signed(((2'd2)));
  assign y4 = (|(4'd2 * (p0?a2:a1)));
  assign y5 = (-5'sd11);
  assign y6 = (3'd2);
  assign y7 = ((4'd5)<=(3'sd2));
  assign y8 = (~|($signed((!p6))?(p3?p14:a2):(+(p1/p15))));
  assign y9 = {3{(+(-2'sd0))}};
  assign y10 = {$signed(p11),(a1),{p15,p5}};
  assign y11 = (-3'sd2);
  assign y12 = {1{($signed(({{a3,a0},(b4+a1)}!==((b0<<<b2)<<(b5>=a0))))>={3{(p13?a3:p16)}})}};
  assign y13 = {4{{1{(p7)}}}};
  assign y14 = ({(b2!==a1)}>>{4{p2}});
  assign y15 = $signed(($signed($unsigned((~|(-(p12?p4:p2)))))));
  assign y16 = (3'd1);
  assign y17 = ((|(({p2,a3}<=$signed(b0))))-(~^{4{b5}}));
endmodule
