module expression_00656(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~&((-2'sd1)<=(4'sd1)))!==(|(~^(5'sd13))));
  localparam [4:0] p1 = ((((2'sd0)<(2'd2))+((2'sd0)>>>(-5'sd11)))>>(((5'sd13)<=(2'd3))>(!(5'd11))));
  localparam [5:0] p2 = ((((^(2'd0))+((4'sd1)==(5'd24)))>(((2'd3)||(2'sd1))^(+(4'd7))))>=((|(|((-3'sd2)-(4'sd1))))>(((2'sd0)!=(-2'sd1))<=((-2'sd1)>>(3'sd1)))));
  localparam signed [3:0] p3 = ((((2'd1)?(3'sd3):(3'sd0))<<((5'd4)?(3'd5):(3'sd3)))&&(-2'sd0));
  localparam signed [4:0] p4 = (~^(!(-(+(^(~&(|((!(3'd1))-(&(-3'sd0))))))))));
  localparam signed [5:0] p5 = (^{1{{1{(+{4{(~((5'd22)?(5'd8):(3'd0)))}})}}}});
  localparam [3:0] p6 = (-2'sd1);
  localparam [4:0] p7 = ((4'd9)>=(3'd5));
  localparam [5:0] p8 = (+((|(-4'sd0))-(-3'sd3)));
  localparam signed [3:0] p9 = ((((3'd6)===(5'sd6))||((-5'sd12)%(2'd1)))>>(((-2'sd0)>>>(-3'sd0))<=((5'sd13)!=(5'd22))));
  localparam signed [4:0] p10 = {2{{1{(4'd7)}}}};
  localparam signed [5:0] p11 = (((-5'sd4)-(-4'sd2))==(!{(3'd6),(4'sd6)}));
  localparam [3:0] p12 = (-{(~^(((-4'sd3)>>(4'd4))===((4'd5)>=(-2'sd0))))});
  localparam [4:0] p13 = ({4{(-3'sd2)}}?((5'sd14)?(2'd3):(-5'sd2)):(4'sd4));
  localparam [5:0] p14 = (+((~&(~^(((3'sd3)||(4'd9))<=(-2'sd1))))&&((~&((3'd5)-(-3'sd2)))/(4'sd2))));
  localparam signed [3:0] p15 = ((4'd0)?(3'sd0):(2'd3));
  localparam signed [4:0] p16 = {1{({1{((4'd0)<=(5'sd6))}}===(((4'sd5)<<(3'd3))===((5'sd10)&&(-3'sd2))))}};
  localparam signed [5:0] p17 = ({(4'd15),(5'd16)}?((-4'sd3)>(5'd6)):{(3'd6),(-5'sd1)});

  assign y0 = ((|(p14>p5))*(|(-p15)));
  assign y1 = ({(|{p13,p4}),(~^(p0<b0)),(a5||p14)}||((!(p14?a0:b5))?(b5-b5):(p14&&p7)));
  assign y2 = (~^(-b4));
  assign y3 = (+(a4<p11));
  assign y4 = (~&($unsigned({(~(p16)),(&(~|p4)),(p15^b0)})==(5'd2 * (~$unsigned(p14)))));
  assign y5 = (-2'sd0);
  assign y6 = {{4{a2}}};
  assign y7 = {4{(2'sd0)}};
  assign y8 = {{(~(|a1)),(~&(~^a4))},{(~|b3),(-a4),{p15,p9}},(~&(!{a1,p17,p12}))};
  assign y9 = (&((p6!=b3)&&(p4)));
  assign y10 = (-2'sd0);
  assign y11 = {2{(b3^b5)}};
  assign y12 = (~&(((~^(-a5))?{(b5+p16)}:(p14-b0))|(~^{(p4?b0:a2),{(~&b3),{b1,a0,b4}}})));
  assign y13 = {{{{{(a5+a0),{{a2}}}}}}};
  assign y14 = (~&(((|(&b4))+(+(-a4)))==((~&(-b5))+(-(a1>b0)))));
  assign y15 = ({{b5,b0,a3}}<<<(a1?a4:a4));
  assign y16 = (((a4-a3)?{b1,b0}:(p16&a2))?($unsigned((&p7))>=(p14<=b0)):{(^a3),{p14,b4},{a3}});
  assign y17 = (b5!=a1);
endmodule
