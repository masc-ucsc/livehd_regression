module expression_00189(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((4'd8)|(2'sd1));
  localparam [4:0] p1 = (5'sd8);
  localparam [5:0] p2 = ((-4'sd3)<<<(5'd11));
  localparam signed [3:0] p3 = (((3'sd1)?(5'd3):(5'd5))?((4'd4)||(4'sd0)):((3'd7)?(2'sd1):(4'd0)));
  localparam signed [4:0] p4 = (-4'sd7);
  localparam signed [5:0] p5 = (~|(5'd2 * (|((3'd5)>(4'd4)))));
  localparam [3:0] p6 = ((4'd4)^~(4'sd5));
  localparam [4:0] p7 = {((3'd6)<(3'd2)),{(-5'sd0),(2'd3)}};
  localparam [5:0] p8 = {(((5'sd10)<<(-2'sd0))<<<(-3'sd0))};
  localparam signed [3:0] p9 = ((|(4'd3))<((4'sd0)?(-2'sd1):(-4'sd7)));
  localparam signed [4:0] p10 = (~|(~^(~&(((6'd2 * (3'd2))>{4{(2'sd0)}})<<<(~&(~|{2{(5'sd1)}}))))));
  localparam signed [5:0] p11 = ((((5'd28)<(4'd6))<((-5'sd2)&(4'sd1)))&&(((2'd2)^(2'sd1))<=((3'd0)|(2'd0))));
  localparam [3:0] p12 = ({4{(2'd3)}}<<<(~|(5'sd12)));
  localparam [4:0] p13 = {{3{{((2'd1)<<(4'sd7)),((-2'sd0)<=(-5'sd10))}}}};
  localparam [5:0] p14 = (-(!(-(((4'd4)?(2'sd0):(-4'sd1))-((-2'sd1)?(-3'sd3):(-5'sd4))))));
  localparam signed [3:0] p15 = {1{((5'sd9)<<<(-3'sd3))}};
  localparam signed [4:0] p16 = (((~|(2'd2))||{(-3'sd0),(5'sd5)})<{((-2'sd0)==(2'd1))});
  localparam signed [5:0] p17 = (-3'sd1);

  assign y0 = $signed($unsigned((($unsigned($signed((p0+p8)))&((a1&&p11)^~(p6|p8)))<=(&$unsigned((&((p14+b3)||(p10<<p5))))))));
  assign y1 = (4'sd7);
  assign y2 = (&$signed((({a2,b1,a4}+($unsigned(a5)<<{a0,b2,b3}))!=={{(+(b2))},(a2?b3:a5)})));
  assign y3 = {{a2,b4}};
  assign y4 = ((+(b4?b0:b5))?{(!(b4?p16:a2))}:{(|(p0?b3:p12))});
  assign y5 = (((b1-b3)<<(b3!=b4))===((a3!=b1)!==(4'd9)));
  assign y6 = (~^(~|((-3'sd2)>=(^((3'sd2))))));
  assign y7 = (2'd3);
  assign y8 = (+((b3?p1:p10)?(b2?p1:p17):(-p8)));
  assign y9 = (5'd1);
  assign y10 = (^{3{(a4>b5)}});
  assign y11 = {(&((|(^(p6|p1)))+({b2,p2,b5}|(p14?b5:p4))))};
  assign y12 = (((p5/a1)?(p8%p3):(a5||p14))^((p3>>a4)>>(a2!=a4)));
  assign y13 = (!(-(((b2&p17)<(p0?p5:p6))?({b1}<={3{p0}}):(+(~(b4+a4))))));
  assign y14 = ({4{(&p17)}}!={3{{p11,p4}}});
  assign y15 = (!((~|((|(a3!==a5))!=((6'd2 * p13)<=(~|b0))))<=({4{b1}}^({4{b2}}+(b0|p11)))));
  assign y16 = (b4?b2:b2);
  assign y17 = (&(!(+(^{2{{(-(+{4{p15}}))}}}))));
endmodule
