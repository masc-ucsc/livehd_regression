module expression_00142(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd7)<<<(3'd7))|{(~(5'd3))});
  localparam [4:0] p1 = (-((3'd6)&((~(2'sd0))+((5'd13)&&(-4'sd3)))));
  localparam [5:0] p2 = (!(-5'sd8));
  localparam signed [3:0] p3 = (((+(|(4'd13)))<=(~^((4'sd2)<(2'd3))))<<(((4'd11)*(-4'sd4))<<<((5'd16)^(4'd3))));
  localparam signed [4:0] p4 = (&(((5'd21)<<<(4'd11))&((4'sd5)?(5'd19):(-5'sd5))));
  localparam signed [5:0] p5 = (((4'd14)<(4'd10))>((2'd0)==(5'd14)));
  localparam [3:0] p6 = (((2'd3)>>(4'd15))?((5'd28)!==(4'sd7)):((-3'sd3)||(3'sd1)));
  localparam [4:0] p7 = (-4'sd1);
  localparam [5:0] p8 = (((2'sd1)===(3'd7))-((-5'sd3)>>>(-5'sd15)));
  localparam signed [3:0] p9 = (~^(({1{{(4'd4),(2'sd1),(2'd3)}}}||((3'd1)&&(-3'sd0)))|(&{4{((2'd1)!==(2'sd0))}})));
  localparam signed [4:0] p10 = ((~({3{(3'sd1)}}<<<((5'sd4)?(3'd5):(-2'sd0))))>>>{4{{4{(-2'sd1)}}}});
  localparam signed [5:0] p11 = ({2{{2{{(3'd6),(-5'sd10)}}}}}<<((((4'd9)<<(2'd1))==={(3'd6),(5'd0),(5'd10)})<<((5'd0)?(2'd1):(-5'sd2))));
  localparam [3:0] p12 = {2{(((4'sd0)?(5'sd9):(2'sd1))<<{2{(3'sd3)}})}};
  localparam [4:0] p13 = (({2{(3'd1)}}^~((4'd10)!=(-3'sd3)))===(~&(!{4{(4'd5)}})));
  localparam [5:0] p14 = (3'd7);
  localparam signed [3:0] p15 = ((&(5'd14))!=={(~&(5'd14)),((-3'sd2)+(3'd5))});
  localparam signed [4:0] p16 = (((~^(|(5'd7)))>=(~|((4'sd1)==(4'd6))))&&(!(~&((~|(3'sd1))>>>(~&(3'd7))))));
  localparam signed [5:0] p17 = {((3'd4)!==(4'd1)),((-3'sd2)?(4'd15):(5'sd7)),((5'd17)^~(4'sd5))};

  assign y0 = {(~(({4{p14}}^~(p15<<<p13))>={3{p7}})),(4'd2 * (p12>p2))};
  assign y1 = {(|(!{{p9,b3},(4'd8)}))};
  assign y2 = (-5'sd4);
  assign y3 = (((a4?b3:b1)>=(~|a5))?{2{{1{b3}}}}:(~^(5'd2 * (b2?b1:a1))));
  assign y4 = {4{b4}};
  assign y5 = (^$unsigned(($signed({b0,a1,a0}))));
  assign y6 = (4'd2 * p2);
  assign y7 = (($unsigned(p2)&&(p13?b5:p0))||((p3?p2:p14)));
  assign y8 = (|(&(~(~^{2{{3{b1}}}}))));
  assign y9 = (($unsigned((-b4)))<<(-(p3*p13)));
  assign y10 = {$unsigned($signed(($unsigned(p9)))),$unsigned(((p14+a3)<(p0<<<p16))),({b4,a1,b4}!==(b5>>a3))};
  assign y11 = (~^$unsigned($signed(($unsigned((+(6'd2 * (b0^a0))))))));
  assign y12 = (-3'sd2);
  assign y13 = (($unsigned($unsigned(a4))-{4{b4}})&&{2{{2{b0}}}});
  assign y14 = (2'd0);
  assign y15 = ({p15}?(-a4):(!b1));
  assign y16 = {1{((&({4{{1{a3}}}}+$unsigned({4{(a4==a4)}}))))}};
  assign y17 = (b1<<p11);
endmodule
