module expression_00354(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd9)!==(-4'sd1));
  localparam [4:0] p1 = {({4{(4'sd1)}}>=(((3'sd3)&(5'd24))-((-2'sd0)===(5'sd14))))};
  localparam [5:0] p2 = {1{{(-5'sd3)}}};
  localparam signed [3:0] p3 = (5'd22);
  localparam signed [4:0] p4 = ((~(~&(4'sd1)))>((((4'd11)>>>(-2'sd1))<<<(&(4'd4)))<=((~|(-2'sd0))*((5'd25)^(2'd3)))));
  localparam signed [5:0] p5 = (-2'sd0);
  localparam [3:0] p6 = ({3{{(2'd2),(2'd0)}}}>>({(+(4'sd5))}>=((5'd21)==(4'd15))));
  localparam [4:0] p7 = (!(3'sd2));
  localparam [5:0] p8 = (~^((-2'sd0)|(5'd18)));
  localparam signed [3:0] p9 = (((3'd5)?(5'd23):(2'd3))?((-4'sd3)?(4'sd3):(5'sd5)):((4'd4)?(2'd3):(-5'sd13)));
  localparam signed [4:0] p10 = ((3'd0)?(2'd1):(-2'sd1));
  localparam signed [5:0] p11 = (((4'sd1)<=(4'd11))/(5'd29));
  localparam [3:0] p12 = (-(({(3'd1),(2'd3)}<<{(5'd17),(4'd10),(5'd10)})^~(3'd0)));
  localparam [4:0] p13 = ((3'd0)>>(5'sd10));
  localparam [5:0] p14 = (|(((~^(-5'sd7))!=(^(2'd2)))=={(-(-5'sd11)),((-5'sd14)^~(3'd1))}));
  localparam signed [3:0] p15 = ((-4'sd3)<<<(5'sd1));
  localparam signed [4:0] p16 = {((&((4'd4)-(3'sd3)))!=(!{(-4'sd1),(-3'sd2)}))};
  localparam signed [5:0] p17 = {1{{(2'd2),(-5'sd11),(5'd0)}}};

  assign y0 = ((b4&&a0)^~(b3<<<b5));
  assign y1 = (2'd0);
  assign y2 = {(5'd10)};
  assign y3 = {({a4,a0}>>>{p13,p6,p14}),((p5?b1:p15)^~(b4<<<p5)),((p8?p9:p2)=={p2,b5})};
  assign y4 = ((p10?a4:b4)&$signed(b3));
  assign y5 = {2{(-((p0^~p13)?(4'd2 * p12):(2'd1)))}};
  assign y6 = (4'd1);
  assign y7 = (|$unsigned($unsigned(((~&{1{{b5,a2,a3}}})))));
  assign y8 = (((p12||p9)-(p4&a3))&&((b5===a2)!=(p8==b1)));
  assign y9 = ((2'd3)&&(b2?p13:p2));
  assign y10 = {{(~&{((~&p5)+{p9})}),{{3{p3}},(p11!=p11),{2{a4}}}}};
  assign y11 = (~(((b1^~a1)?(-(~&a0)):(4'd2 * a0))!==(^(($unsigned(b5))?(&(a1?b0:a2)):(b0!=a2)))));
  assign y12 = (~^(+({2{(b2>>a5)}}|(|{1{(a5?a0:b2)}}))));
  assign y13 = {{2{{1{{{1{{a1}}},(b5<a4),{4{a0}}}}}}}};
  assign y14 = (!(p11%a1));
  assign y15 = (~|((&(((-$unsigned((~|$signed((~&(+$signed($unsigned((~^((~&((~&p3))))))))))))))))));
  assign y16 = (!((+(p15|b5))==(-(-a0))));
  assign y17 = ((a4?a1:a2)|(2'd1));
endmodule
