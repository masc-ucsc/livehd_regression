module expression_00732(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd9)|(3'sd1))%(-5'sd0));
  localparam [4:0] p1 = (((5'sd15)&(-5'sd12))>>((4'd12)^~(-5'sd7)));
  localparam [5:0] p2 = {{{(4'sd5),(-2'sd0),(4'd14)},{(4'sd3),(3'd5),(3'd0)}},(4'd9),{(-(4'sd1)),(4'sd0)}};
  localparam signed [3:0] p3 = (4'd2 * {1{(2'd2)}});
  localparam signed [4:0] p4 = (((-2'sd1)?(4'd6):(3'sd2))?(~|(-2'sd1)):(~^(5'sd9)));
  localparam signed [5:0] p5 = ((((-5'sd11)?(5'd1):(4'd6))?{3{(3'd3)}}:((5'd28)!==(4'd11)))+(((4'd13)|(-5'sd4))<=((-3'sd2)!==(5'd12))));
  localparam [3:0] p6 = ((!((|(5'd30))^((-3'sd0)^~(2'd1))))^~(((4'sd6)>(-2'sd0))>>(~&(~|(5'sd2)))));
  localparam [4:0] p7 = (|(((2'd0)?(2'sd0):(2'd1))/(-3'sd2)));
  localparam [5:0] p8 = (|(((^(-3'sd3))?{1{(2'd2)}}:{1{(-4'sd7)}})<<<(~|(3'd3))));
  localparam signed [3:0] p9 = (|{{(&{(4'd1),(2'sd0),(5'sd4)}),{2{{3{(3'd7)}}}}}});
  localparam signed [4:0] p10 = {(5'd0),(-4'sd2),(-2'sd0)};
  localparam signed [5:0] p11 = (-5'sd7);
  localparam [3:0] p12 = ((4'd2 * ((3'd1)?(4'd5):(2'd3)))||(((3'd6)<<<(3'd0))!==((2'd3)?(2'sd0):(3'sd1))));
  localparam [4:0] p13 = (!(~^(3'sd1)));
  localparam [5:0] p14 = (~&((4'd2 * (+((5'd9)?(3'd4):(2'd1))))?(((2'd2)&&(4'sd0))?(+(5'sd10)):((3'sd3)?(-5'sd0):(5'd3))):(~^(~|((5'd6)?(5'd10):(4'd5))))));
  localparam signed [3:0] p15 = ((+((!(3'sd3))<=((-5'sd4)<<<(3'sd1))))?(((3'd5)^(5'd19))-((4'd15)==(4'd0))):((3'd2)/(4'sd3)));
  localparam signed [4:0] p16 = ((((5'd9)<<(-3'sd3))==(~^(-2'sd1)))>>{((5'd29)|(4'sd3)),((-2'sd0)<<<(5'd14)),((-2'sd1)?(5'd7):(5'sd3))});
  localparam signed [5:0] p17 = {(~|{3{{2{((2'sd1)>(5'd1))}}}})};

  assign y0 = $unsigned(((b1==b4)));
  assign y1 = ({1{(+((a0<<<p6)<<{3{b4}}))}}<<<{(p11||p1),{1{p15}},(3'sd2)});
  assign y2 = (5'd23);
  assign y3 = $unsigned({1{((p13>p14)||(p14^p2))}});
  assign y4 = {$signed(((p7-a5)&$unsigned((p17<p2))))};
  assign y5 = (6'd2 * b2);
  assign y6 = (^{1{({4{p8}}>>>(-p14))}});
  assign y7 = (+(~{(((b2<<<p9))<<((p7^p11))),({p14,p8,p10}<<{p5,p8}),(|(4'd2 * $unsigned($signed(p10))))}));
  assign y8 = (&b3);
  assign y9 = {(((a5&&b0)-(~^(b5>b5)))>>>((b3===b2)||(a5-a2)))};
  assign y10 = {((b2&&b5)!==(b5===b1)),((a4==p14)<(3'd1))};
  assign y11 = ((4'd2 * p7)!=(p7^~p9));
  assign y12 = ((-((^(a3?a3:p10))<={4{p1}})));
  assign y13 = (b5?a0:a3);
  assign y14 = ((+b3)+(-4'sd2));
  assign y15 = (3'sd1);
  assign y16 = {{(4'd7)},{1{(~^p0)}},{4{a3}}};
  assign y17 = ((({a2}<={a2,a2})<<(~^{b2,b4,b1}))&{(|(~^{(+b1),(b4+a0)}))});
endmodule
