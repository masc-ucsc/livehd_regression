module expression_00689(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({1{((5'd15)?(3'sd3):(3'd5))}}?({2{(-3'sd0)}}!==((-2'sd1)?(4'd14):(-4'sd3))):(2'd1));
  localparam [4:0] p1 = (+((-5'sd13)?(^((4'd6)?(5'd30):(4'sd3))):((3'd3)?(2'sd1):(-2'sd1))));
  localparam [5:0] p2 = ((4'd11)>(3'd2));
  localparam signed [3:0] p3 = ((4'd11)?((~^(3'sd1))|((5'sd0)>>(5'sd4))):(-5'sd15));
  localparam signed [4:0] p4 = {({{(4'd0),(-3'sd0),(-5'sd7)}}|((&(3'd6))-((2'd3)===(3'd1))))};
  localparam signed [5:0] p5 = ({(3'sd2),(3'sd2),(-5'sd8)}||((2'sd0)?(2'd2):(2'sd1)));
  localparam [3:0] p6 = {{3{({4{(-5'sd6)}}&&((5'd9)>=(2'd0)))}}};
  localparam [4:0] p7 = (2'sd1);
  localparam [5:0] p8 = {4{{1{(5'sd1)}}}};
  localparam signed [3:0] p9 = {{(((2'd3)?(2'sd0):(2'd3))!==((3'd4)>(5'sd7)))},{((-3'sd0)?(4'd14):(4'd8))}};
  localparam signed [4:0] p10 = {((-3'sd0)?(^(4'd5)):((5'd19)>(5'sd3))),({(4'd6),(4'd10),(2'd3)}<<(~|(|(3'd6))))};
  localparam signed [5:0] p11 = ({(-5'sd14),(3'd7)}<=(2'd2));
  localparam [3:0] p12 = ((3'd0)<<<(5'sd10));
  localparam [4:0] p13 = (3'd4);
  localparam [5:0] p14 = (6'd2 * (~&{4{(4'd2)}}));
  localparam signed [3:0] p15 = {1{((5'sd7)||(3'd0))}};
  localparam signed [4:0] p16 = ((4'd2 * (3'd1))?(~(4'd4)):{(5'd31)});
  localparam signed [5:0] p17 = {{(-4'sd2)},(+(-2'sd0)),(-(4'd9))};

  assign y0 = $signed((5'd14));
  assign y1 = ((5'd2 * (b1*a0))^~$signed((!$signed(b0))));
  assign y2 = (^({2{{4{p9}}}}<<<((a2>>>b5)===(^(b1+b3)))));
  assign y3 = (~^(&(({p0,p8,a0}?(+a1):(a3^~b2))>=($signed(a1)?{p8,a0,a4}:(b1?p9:b0)))));
  assign y4 = (~^(+(&(^(!({1{({3{a4}}!=={2{b0}})}}||(+(~^{4{a3}}))))))));
  assign y5 = (|{2{({(^a3)}&(b1+p1))}});
  assign y6 = (!(!(($unsigned(p4)|(-3'sd3))?(~(-$signed(a2))):($signed((b3))))));
  assign y7 = ({1{{4{(p10^p11)}}}}+{1{{1{((p7^p8)<<<{4{p0}})}}}});
  assign y8 = {3{((^(~|a5))>=(b1===b4))}};
  assign y9 = {3{(|(-4'sd6))}};
  assign y10 = {2{((p14?p17:b4)&&{3{p8}})}};
  assign y11 = ((-3'sd3)?(5'sd2):(b0?p2:a4));
  assign y12 = (a3<<b4);
  assign y13 = (3'd1);
  assign y14 = ({2{{4{b4}}}}<((((b4<<p5))?(^{2{b2}}):(b2<p12))));
  assign y15 = (4'd2 * (a1?b2:a2));
  assign y16 = {3{((a2==b0)!==(a1|b0))}};
  assign y17 = (^(~&({2{(|b3)}}?(!(+(p4?a5:b1))):{4{a4}})));
endmodule
