module expression_00045(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((5'sd14)-(-5'sd7))?((5'd13)?(2'd0):(2'd1)):((4'd3)?(4'd2):(5'sd12)))?(6'd2 * ((2'd1)?(2'd2):(2'd0))):(((4'sd4)%(5'd11))&&((2'd1)>>>(-3'sd1))));
  localparam [4:0] p1 = (~|(~^(&{1{{2{(~^(5'd23))}}}})));
  localparam [5:0] p2 = (&{(~(+(((!(3'd5))^~{(2'd0),(5'd11)})<<<((~(4'd5))==((3'd6)!==(-2'sd1))))))});
  localparam signed [3:0] p3 = {4{{(3'd2),(-2'sd1),(-3'sd0)}}};
  localparam signed [4:0] p4 = (4'd5);
  localparam signed [5:0] p5 = ((~|(4'sd4))!==((5'sd13)<<<(3'd3)));
  localparam [3:0] p6 = {1{((~(^(-3'sd3)))?{3{(-5'sd8)}}:{3{(-5'sd15)}})}};
  localparam [4:0] p7 = ((((-2'sd0)?(4'sd4):(5'd2))==(-3'sd1))^~((2'sd0)?(-2'sd0):(4'd13)));
  localparam [5:0] p8 = {3{{(-3'sd0),(3'd7)}}};
  localparam signed [3:0] p9 = (&((2'd0)>>(4'sd3)));
  localparam signed [4:0] p10 = (-{1{({(5'sd4),(5'd5)}?((2'sd1)?(2'd0):(3'd6)):{4{(-3'sd0)}})}});
  localparam signed [5:0] p11 = (5'sd10);
  localparam [3:0] p12 = {{{(~^(5'd31)),(&(4'd1)),{(5'sd7),(-5'sd9)}}},(!{{(|(4'sd0)),(~|(4'sd0)),{(5'd31),(-4'sd1),(-5'sd6)}}})};
  localparam [4:0] p13 = (((2'd0)!==(4'd8))==={(5'd2),(5'sd14)});
  localparam [5:0] p14 = {4{(3'sd1)}};
  localparam signed [3:0] p15 = (~(~^{(-3'sd1),(4'd15),(5'sd9)}));
  localparam signed [4:0] p16 = {4{(2'd2)}};
  localparam signed [5:0] p17 = {4{(3'd6)}};

  assign y0 = ({2{(a2|b1)}}^~({4{a4}}?(~|a4):(|b3)));
  assign y1 = ({(a4?b5:b2),(p3?a2:a3),{p16,b1,b1}}?((a5)?(a1?a5:a1):{p16}):$unsigned($unsigned({a4,a1,b3})));
  assign y2 = (((!(^b3))?(&(b5?b4:a2)):(|(|a3)))+(|((+(~(!p12)))==(|(~&{a5,a3,a4})))));
  assign y3 = (((~b0)?{b3,a5,b1}:{4{a0}})?{(p7?b4:p12),(~&p15),{2{p8}}}:{3{(a0?p16:p10)}});
  assign y4 = (!({p3}?{a5}:(p8>=p2)));
  assign y5 = (((p14?p6:p5)?(p16?b3:b1):(a5?a0:b3))?{4{(p2?p3:a1)}}:{2{{2{a3}}}});
  assign y6 = ((a2%p4)==(&(5'd4)));
  assign y7 = ({((p16?p5:b0)?{4{p6}}:(p11?p2:b5))}^((|{1{(~&p14)}})^(~{1{(-5'sd14)}})));
  assign y8 = {1{({1{(~^p16)}}>>>(a2<=a2))}};
  assign y9 = (((^p16)>>(p1<a1))?((b0?b2:p10)>>{4{p12}}):{4{p10}});
  assign y10 = (p12||a3);
  assign y11 = $signed($signed({2{(&{4{p0}})}}));
  assign y12 = $signed((((b0?p12:p10)||(|{p8,p10,a5}))?{(p14>=p12),{1{{p5,a5}}}}:(^({4{p9}}?{4{p5}}:(p0)))));
  assign y13 = {{(~&a0),{4{p2}},{b5,a0,p16}},(~&{3{p14}})};
  assign y14 = ((5'd18));
  assign y15 = {4{(3'd2)}};
  assign y16 = (+((^(4'sd7))));
  assign y17 = ((5'd2 * (5'd2 * p13))^{(p17+p9),(p13>>p16),$unsigned((p17^p17))});
endmodule
