module expression_00487(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-2'sd1);
  localparam [4:0] p1 = (~^(((~|(5'd26))?(-(3'sd1)):((-3'sd1)<(5'sd12)))|{(|(4'd5)),((4'sd7)>>(3'sd2)),(~|(2'd3))}));
  localparam [5:0] p2 = (5'd13);
  localparam signed [3:0] p3 = {(~&((3'd2)===(4'd2)))};
  localparam signed [4:0] p4 = {({2{(3'd4)}}<<<{3{(4'sd1)}})};
  localparam signed [5:0] p5 = (5'd2 * ((2'd0)?(3'd2):(2'd2)));
  localparam [3:0] p6 = ({4{{(2'd3)}}}&{4{((-5'sd15)?(5'd26):(4'd6))}});
  localparam [4:0] p7 = (+((2'sd1)>>(((3'd6)?(2'sd1):(5'sd6))<<<(^(~|(-4'sd5))))));
  localparam [5:0] p8 = ((-3'sd1)?(2'd2):(-4'sd4));
  localparam signed [3:0] p9 = (~&{((-(2'd2))>>>((5'sd4)===(4'd11))),((3'sd2)?(4'sd0):(5'd26)),{3{(2'sd1)}}});
  localparam signed [4:0] p10 = ((~((3'd4)|(3'd3)))&&(&(-{(3'd1),(3'd7),(4'd1)})));
  localparam signed [5:0] p11 = {1{(({((3'd4)+(-5'sd14))}^{4{(2'd0)}})>((4'd2 * (3'd7))<<((3'sd3)==(5'd23))))}};
  localparam [3:0] p12 = (((5'sd11)<=(5'sd0))==={4{(-4'sd5)}});
  localparam [4:0] p13 = (((2'sd0)<=(-5'sd1))*((3'd6)/(5'd15)));
  localparam [5:0] p14 = (((2'd1)?(2'd2):(2'sd1))?(-4'sd0):(~&((5'd28)||(4'd6))));
  localparam signed [3:0] p15 = {((2'sd1)?(-2'sd1):(5'sd0)),((5'sd4)?(2'sd1):(3'd4)),((4'sd4)&(-3'sd3))};
  localparam signed [4:0] p16 = ((5'd15)!==(-(((5'd7)>>(4'sd6))>(~|{2{(-2'sd1)}}))));
  localparam signed [5:0] p17 = (((!(4'd14))?((-2'sd0)===(2'd1)):{(3'd3),(2'sd1)})|{(~^((2'd1)!=(4'sd3))),(^{(3'd2)})});

  assign y0 = (a3&p16);
  assign y1 = (({3{b5}}<<{3{b2}})==={{3{{2{a0}}}}});
  assign y2 = ((p5||p12)|(p3>a4));
  assign y3 = {1{({3{{4{b4}}}})}};
  assign y4 = {{p13,p3,a3}};
  assign y5 = (4'd2 * (b1<<a2));
  assign y6 = (5'sd10);
  assign y7 = (3'd6);
  assign y8 = ((a0<b1)==(p17^a4));
  assign y9 = ((5'd20)<<<{4{p16}});
  assign y10 = ((((&b3)=={b4,a1,a5})&&{$signed(a2),(~|b3)})!={1{(~(~|((a0+b1)<={1{a3}})))}});
  assign y11 = (3'd2);
  assign y12 = (({b1,b3,b2}<<<(!(~|(~|a2))))===(!(~&((!{3{a4}})<={b1,b3,a4}))));
  assign y13 = ((b0!=a4)<=(p7==p3));
  assign y14 = {4{((a4>a4)||(p4^b0))}};
  assign y15 = (~|(4'd4));
  assign y16 = (p16|p4);
  assign y17 = ((p0>=p16)?(a0>=p13):(p16?p4:p12));
endmodule
