module expression_00959(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{(-4'sd5)}};
  localparam [4:0] p1 = ((((2'sd0)<=(-4'sd6))>=(~^(5'd12)))!==(((-5'sd0)>(4'sd3))|(&(4'sd4))));
  localparam [5:0] p2 = (4'sd3);
  localparam signed [3:0] p3 = (((5'd7)!==(-3'sd2))?((-3'sd1)>>(-4'sd6)):{(3'd5),(-4'sd5)});
  localparam signed [4:0] p4 = (((-4'sd4)>=(2'sd1))/(-2'sd1));
  localparam signed [5:0] p5 = (((5'sd6)^~(3'd2))!==(3'sd2));
  localparam [3:0] p6 = {((5'd8)||(-(~(2'd2))))};
  localparam [4:0] p7 = (((4'd2 * (4'd8))<(~&(-2'sd1)))>(^(~((2'sd1)>(2'sd0)))));
  localparam [5:0] p8 = (-(~&((2'd2)-((2'd2)||(-2'sd1)))));
  localparam signed [3:0] p9 = {({((3'sd3)|(5'sd3))}<<{(4'd5),(5'sd6),(-2'sd1)})};
  localparam signed [4:0] p10 = {(4'd10)};
  localparam signed [5:0] p11 = (((-5'sd0)-(2'sd1))+((2'd2)||(4'd3)));
  localparam [3:0] p12 = (~|((3'sd0)?(-4'sd4):(-2'sd1)));
  localparam [4:0] p13 = (((3'sd3)<=(-5'sd2))%(-4'sd1));
  localparam [5:0] p14 = {((3'd1)?(4'sd0):(3'd7)),{{(-5'sd8),(4'd0)}},(2'sd1)};
  localparam signed [3:0] p15 = (~&((((-5'sd12)!=(2'd3))|(5'sd8))?(~^((-3'sd0)?(4'd13):(4'd1))):(2'sd1)));
  localparam signed [4:0] p16 = ((~^((4'd9)||(-3'sd3)))>>((-3'sd3)>>>(4'd14)));
  localparam signed [5:0] p17 = {2{(-3'sd0)}};

  assign y0 = {3{{3{a4}}}};
  assign y1 = {4{({1{p4}}<=(2'd1))}};
  assign y2 = (~^{(|(^(~|$unsigned(a3)))),((~(p2<b2)))});
  assign y3 = ((~|(p8?p7:p6))>>((3'd5)&&(p10==p10)));
  assign y4 = (&p5);
  assign y5 = ((5'd2 * (p1!=p12))?((b0!=b1)?(a0+a1):(p9|b4)):($unsigned(b2)*(p10*p17)));
  assign y6 = (~&($signed((~^b3))?$unsigned($unsigned(p15)):(~|(p4?a2:p13))));
  assign y7 = {1{{4{((a1>b4)==={a0,b3})}}}};
  assign y8 = ((^((&(a3!=a5))>=(p10^~b1)))<<((b3<a1)>(p5+a3)));
  assign y9 = {((&(~|(-p16)))),((~|p6)<=(p10>p17)),{3{{3{p2}}}}};
  assign y10 = ({4{(a5)}}?($signed({1{p15}})<<<(p15!=p12)):$signed({3{(^b1)}}));
  assign y11 = (5'd19);
  assign y12 = (-(~^(^((p13*a2)*(p11?b0:p8)))));
  assign y13 = (-4'sd1);
  assign y14 = $unsigned(p7);
  assign y15 = (+(~&(+(3'd1))));
  assign y16 = (((~|(|(-(p5/p12))))|((p10+b5)/p11))+(((b4>>>a2)%b2)>>>((~&b0)<(&b0))));
  assign y17 = ((a0?b0:p7)?$unsigned((a3>a0)):((b1>=p11)!=(b4)));
endmodule
