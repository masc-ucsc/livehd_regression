module expression_00115(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(~&((-((3'd4)==(4'd14)))%(4'sd4))));
  localparam [4:0] p1 = (|(+(!({{(3'd6),(2'sd0)},(~|(4'd11)),{(4'd0),(4'd11),(-4'sd6)}}=={{(+(4'sd1)),{(5'd16),(5'sd6),(5'd11)}}}))));
  localparam [5:0] p2 = ((-((5'sd12)?(4'd6):(-2'sd1)))>>(((-3'sd2)?(3'd7):(4'd9))?{1{(2'd1)}}:(~|(-4'sd0))));
  localparam signed [3:0] p3 = {2{((2'sd0)?(5'sd2):(5'sd6))}};
  localparam signed [4:0] p4 = {(^((2'd2)||(-3'sd2))),(~^{(5'd18),(4'sd6)})};
  localparam signed [5:0] p5 = (~^(5'd20));
  localparam [3:0] p6 = ((~^(((-3'sd3)<(2'sd1))+(~^(5'sd3))))&&{3{{(3'd5),(3'd5),(3'd4)}}});
  localparam [4:0] p7 = ((~(-2'sd0))!=(+(-4'sd1)));
  localparam [5:0] p8 = {(5'd12),(3'sd1),(3'd7)};
  localparam signed [3:0] p9 = (~&(~|((((-4'sd1)/(-4'sd5))<=(~|((5'd26)&(4'd15))))>=((!(|(4'sd0)))&((-3'sd3)>>(-2'sd1))))));
  localparam signed [4:0] p10 = (+({(5'sd3),(-2'sd0),(3'd2)}=={1{((-5'sd7)-(2'd1))}}));
  localparam signed [5:0] p11 = (5'd2 * ((2'd1)&(3'd1)));
  localparam [3:0] p12 = {4{(-5'sd13)}};
  localparam [4:0] p13 = (2'd3);
  localparam [5:0] p14 = (((2'sd0)%(-4'sd5))*((5'd4)>(5'sd1)));
  localparam signed [3:0] p15 = ({(((5'sd1)<<(-4'sd0))<=((4'd6)<(2'd1)))}^({(2'd1)}?(~&(5'sd12)):((2'd0)!==(4'd12))));
  localparam signed [4:0] p16 = (-2'sd1);
  localparam signed [5:0] p17 = (5'sd9);

  assign y0 = (p12||p0);
  assign y1 = (4'd4);
  assign y2 = ((((p10?p10:a0)^(a5?a2:p1)))||((-(p4?b4:a5))));
  assign y3 = ((((a4?b5:b2)^~(b5<<<b0))&&({a5,p10,a2}-(a4?b1:a3)))^{(+(a2<p14)),(b2||a2),(p11==a4)});
  assign y4 = (((p16?b0:b1)^~(a0?b3:a0))|(6'd2 * $unsigned((b0?p15:a4))));
  assign y5 = (2'd1);
  assign y6 = (+{(~&$signed(p4)),$unsigned({b1,p3}),(|{p2,p1})});
  assign y7 = (((p8?p16:p15)-(p1*p10))?($signed($signed((p9<=p1)))):((p4?p2:b1)?$unsigned(p3):(p13>=p6)));
  assign y8 = ((a0||b1)?(p10>>>p17):(a5!==b2));
  assign y9 = $unsigned(({((-2'sd1)|(a3===b0))}>>>((p1<<a5)&(b0===b0))));
  assign y10 = (((b5+a1))*(b4/b1));
  assign y11 = (+{1{{4{p5}}}});
  assign y12 = ((|(+(-({a1,a2}|(a2|b5)))))===(({b4}<<<(a5>a1))<<({b1,a0}|(b5^b0))));
  assign y13 = ($unsigned($signed((4'sd6)))?(4'sd1):((4'sd1)<=(b4?p15:p3)));
  assign y14 = ((5'd0)<<<(4'd0));
  assign y15 = (({4{p2}}||{2{p10}})>=((b0^p7)&&(a5&a2)));
  assign y16 = ((3'd2)&(|((~|(b5?b3:a4))?(-2'sd1):(a4%a2))));
  assign y17 = {2{{{(~&{a5,p0,p15}),$signed({b2,a3})}}}};
endmodule
