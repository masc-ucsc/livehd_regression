module expression_00936(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(3'd3));
  localparam [4:0] p1 = (4'd2 * (4'd6));
  localparam [5:0] p2 = {{(2'd0),(2'd1)}};
  localparam signed [3:0] p3 = (((5'd21)!==(-4'sd1))?((-5'sd0)?(3'd2):(3'd7)):((2'sd0)?(2'd1):(5'd21)));
  localparam signed [4:0] p4 = ({3{((2'd2)||(3'd4))}}>>(&(^{3{((4'd12)==(4'd1))}})));
  localparam signed [5:0] p5 = ({3{(3'sd2)}}!==(((4'sd5)>>>(4'sd5))||((4'sd5)!==(4'sd3))));
  localparam [3:0] p6 = (~^(|(~&(((4'd15)?(-2'sd1):(5'd27))?(!(-5'sd4)):((3'd3)?(-5'sd4):(-2'sd1))))));
  localparam [4:0] p7 = {{((4'd8)+(2'sd0))},(((3'd4)^(3'd1))|(&(3'sd2)))};
  localparam [5:0] p8 = {(((3'd5)===(3'sd1))<<<{(2'sd0),(5'sd14),(-5'sd2)}),((-(5'd2 * (2'd1)))<<<{(5'd14),(2'd2),(2'd1)})};
  localparam signed [3:0] p9 = {4{(~(+(4'd0)))}};
  localparam signed [4:0] p10 = (((!(4'd6))<=((2'd2)?(-5'sd8):(-3'sd2)))?{(~&(4'd8)),(~(4'd9)),{2{(-3'sd3)}}}:({1{(4'sd1)}}&(|(3'sd3))));
  localparam signed [5:0] p11 = (+(({1{(3'd7)}}!==((-5'sd11)==(-5'sd12)))-(((-3'sd0)===(2'd1))+{3{(4'd5)}})));
  localparam [3:0] p12 = (((2'sd1)^(2'sd1))>(4'sd4));
  localparam [4:0] p13 = {1{{4{((2'sd0)>=(5'sd5))}}}};
  localparam [5:0] p14 = {4{(-2'sd1)}};
  localparam signed [3:0] p15 = (|(|(((~&(5'sd11))<((4'd13)>>(2'sd0)))!=(|(6'd2 * (!(5'd8)))))));
  localparam signed [4:0] p16 = {3{{{(5'd30),(2'sd0)}}}};
  localparam signed [5:0] p17 = ((5'd28)?(2'd2):(5'd14));

  assign y0 = (&(|(($unsigned((|((a1%p0))))<((!(~&p1))|(!(5'd2 * a1)))))));
  assign y1 = ((a5/a5)%b0);
  assign y2 = (~(-5'sd11));
  assign y3 = (-((~|(-$signed((-4'sd6))))<<(2'sd1)));
  assign y4 = {3{b0}};
  assign y5 = ({1{{4{p9}}}}?{(p17?p10:p17)}:(p3>>p9));
  assign y6 = ({p17,p7}==(-b1));
  assign y7 = $signed((p4?a3:b5));
  assign y8 = (^(-({({3{p14}}-{a1,p5,p2})}^~(~^({p11,p0,p10}+(p0<<a1))))));
  assign y9 = (b3>>a1);
  assign y10 = (~&(!(^(-(|(p9>>p11))))));
  assign y11 = ((p16|p16)?(p7==p4):(-p12));
  assign y12 = ((a3<=p2)?(p9<=b1):(b1|p3));
  assign y13 = (~(!(~(&(+(|(~^(~^(~&(+(-p7)))))))))));
  assign y14 = (2'd1);
  assign y15 = (-5'sd11);
  assign y16 = ((~&$signed(a5))>(+(p0>>>b0)));
  assign y17 = $unsigned(((^(~&p5))));
endmodule
