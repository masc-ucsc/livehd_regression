module expression_00859(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&((&(2'd2))<{2{(5'd16)}}));
  localparam [4:0] p1 = ((&(-5'sd1))!==((-2'sd1)-(3'sd1)));
  localparam [5:0] p2 = ((2'd3)?(-4'sd1):(4'sd7));
  localparam signed [3:0] p3 = {({{(3'sd2),(5'd22)}}>>>(&((4'd4)<(3'sd3)))),{{(2'sd0),(5'd17),(-5'sd13)},(|(~|((-4'sd7)!=(5'sd6))))}};
  localparam signed [4:0] p4 = ((4'd6)===(5'sd5));
  localparam signed [5:0] p5 = {({1{((4'd8)===(3'd7))}}?(((5'd27)?(5'sd0):(4'sd3))>>>((2'd0)^~(5'd11))):((4'd10)?(3'sd1):(-2'sd1)))};
  localparam [3:0] p6 = {(((2'd0)+(2'sd0))>>((2'sd0)<<(-3'sd0))),{{(4'd7),(-4'sd4),(-2'sd1)},((3'd3)||(3'd5))},(((5'sd6)?(2'd2):(5'sd9))?((5'd22)?(2'sd0):(5'd21)):{(4'd7),(4'sd5),(4'd5)})};
  localparam [4:0] p7 = ((~^((5'd21)>=(3'd7)))?((4'd8)||(5'd6)):((2'd2)^(5'd25)));
  localparam [5:0] p8 = ((&((~|(~^(-3'sd0)))<<(-(!(5'd27)))))<((~{(4'd11),(2'd0),(3'd7)})<<(^{(4'd7),(2'd0),(2'd2)})));
  localparam signed [3:0] p9 = ((2'd2)^(-2'sd0));
  localparam signed [4:0] p10 = ((~(3'd3))>=((3'd0)?(2'sd0):(3'd1)));
  localparam signed [5:0] p11 = (((~|(5'sd13))>=((3'd6)?(2'sd0):(5'd30)))?(+((3'd5)===(4'd4))):(~((-2'sd1)?(-3'sd1):(4'd4))));
  localparam [3:0] p12 = ((((3'd0)?(-2'sd1):(2'sd0))?((3'd5)||(-4'sd6)):((3'd0)!==(-3'sd3)))<<{1{((~^((3'sd1)?(5'd14):(4'sd2)))<{3{(-5'sd11)}})}});
  localparam [4:0] p13 = (((4'd2)?((4'd8)>>(3'd0)):{4{(-2'sd1)}})==={3{((-2'sd0)^(3'd4))}});
  localparam [5:0] p14 = (2'd1);
  localparam signed [3:0] p15 = {(+((2'd3)^~(-5'sd6))),((2'd3)?(3'sd2):(4'sd2)),(~^{(3'd7),(2'd3)})};
  localparam signed [4:0] p16 = (((4'd10)<(-4'sd4))*((5'd20)-(3'd4)));
  localparam signed [5:0] p17 = (((4'd1)<(5'sd8))>=(4'd6));

  assign y0 = ((b2<a2)>=(b2?p10:p15));
  assign y1 = {1{($unsigned({3{b0}})>>((a3&&a1)>>>(a2||p1)))}};
  assign y2 = ((^(~|(b3&p15)))<<({b2,b3}&&(a4+b3)));
  assign y3 = ((p10?p6:p9)==(p13?p9:a2));
  assign y4 = ((|{{{p6},{a3,p11}},{1{{a1,a4}}}})^~{2{{{a2,p0,p15},(-p7)}}});
  assign y5 = (&{4{(a5?a3:a5)}});
  assign y6 = ({b2,b0}-(b2==a3));
  assign y7 = (-5'sd2);
  assign y8 = (~&(5'sd13));
  assign y9 = {4{(-3'sd2)}};
  assign y10 = (+(|((a4!==b2)-(~^{a3}))));
  assign y11 = ((-4'sd0)!==((a5?a4:a0)?(a2|b1):(b2?b5:b3)));
  assign y12 = ({p5,p2,p13}?{3{p11}}:{3{p11}});
  assign y13 = ((&(&(a0-a2)))?((p6>a1)==(p1?a1:p2)):((p17?p17:b5)>>(p9^~b5)));
  assign y14 = ((-2'sd0)<=((-3'sd1)|(2'd2)));
  assign y15 = $unsigned(((~(+({3{p14}}<<<(b2>>a0))))||(~&(-$signed((6'd2 * $unsigned((p5^p17))))))));
  assign y16 = {(({b4,b4}<=$signed(p4))||(-{(p13),$unsigned(p3)}))};
  assign y17 = {{{p11,b1,b5}},{{b3,p12}},{{p14,p2}}};
endmodule
