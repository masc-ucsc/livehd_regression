module expression_00398(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((~^(~|(4'd7)))+{4{(5'sd0)}})<<<{2{{3{(2'd3)}}}});
  localparam [4:0] p1 = ((~&(&(5'd30)))<<(~^((-4'sd7)?(2'sd1):(-4'sd2))));
  localparam [5:0] p2 = ({{1{(4'd6)}},{(3'd3)}}?{2{((5'd18)<<(2'd2))}}:((-3'sd0)?(4'd4):(5'd1)));
  localparam signed [3:0] p3 = (((5'd31)?(2'd0):(4'd9))!=((5'd16)?(3'd4):(4'd12)));
  localparam signed [4:0] p4 = ({2{{(5'sd7),(5'd6),(-4'sd0)}}}^(~^({(!(2'd0))}-{4{(2'd1)}})));
  localparam signed [5:0] p5 = (5'd14);
  localparam [3:0] p6 = (^{{(2'sd0),(3'sd1),(3'd3)},(~^(2'sd1))});
  localparam [4:0] p7 = {(4'd2 * {(3'd5),(4'd0),(5'd24)})};
  localparam [5:0] p8 = ((((3'd1)?(5'sd6):(3'sd2))?{2{(2'd0)}}:{1{(4'd11)}})+{(((4'sd1)?(-3'sd2):(-4'sd2))?((3'd2)|(-3'sd3)):{4{(-3'sd1)}})});
  localparam signed [3:0] p9 = {4{(2'd1)}};
  localparam signed [4:0] p10 = (~^(~&(5'sd8)));
  localparam signed [5:0] p11 = ((5'd2 * (2'd3))?((5'd31)-(3'd4)):((3'sd3)?(5'd18):(5'd14)));
  localparam [3:0] p12 = {({(5'd1),(2'd2)}-{4{(5'd29)}})};
  localparam [4:0] p13 = {{2{{((4'd6)==(4'd3)),((-2'sd0)>>>(3'sd2))}}}};
  localparam [5:0] p14 = {(4'd7),(-4'sd5),(4'sd2)};
  localparam signed [3:0] p15 = (-2'sd1);
  localparam signed [4:0] p16 = ((6'd2 * ((2'd3)?(5'd27):(4'd12)))?((2'sd0)?(3'd3):(3'd4)):(-3'sd1));
  localparam signed [5:0] p17 = (~&(5'sd2));

  assign y0 = (~&{2{(^(~&((b3?p9:b5)>>{4{b3}})))}});
  assign y1 = (b5?p17:p3);
  assign y2 = (($signed(b3)>(a0===b1))-({4{a5}}|(~|b1)));
  assign y3 = ((b5^a1)>(^(|p3)));
  assign y4 = (~(~|b5));
  assign y5 = (p9?p3:a4);
  assign y6 = (2'd1);
  assign y7 = {3{{2{(p11?p14:b0)}}}};
  assign y8 = (p9?p2:p14);
  assign y9 = {2{{(~p2)}}};
  assign y10 = ($signed(($unsigned({1{a0}})||{4{p13}})));
  assign y11 = ({2{p3}}?{3{p8}}:{4{p2}});
  assign y12 = {b0};
  assign y13 = (!{((~{{b0,p13}})?((~&a2)<=(p2<<a3)):(&(p11?a3:p1)))});
  assign y14 = (~&(-4'sd0));
  assign y15 = ({(a3-b5),(5'd2 * a1)}?(a2?a5:p3):((3'd7)>>(&p9)));
  assign y16 = ({p5}|{3{p0}});
  assign y17 = (|(((p11?p5:a4)?{p16,p14,p4}:(a1||p5))?(&({3{p11}}?(~&p14):{b0})):(5'd2 * (p13!=a1))));
endmodule
