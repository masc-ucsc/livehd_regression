module expression_00054(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({(2'd1),((3'd5)+(4'd2)),(3'd1)}-(((2'd0)^~(3'sd1))>((3'sd3)>>>(-4'sd0))));
  localparam [4:0] p1 = (&(((2'd3)?(2'd3):(2'sd1))?((-2'sd0)?(3'd6):(-3'sd2)):(~|((3'd5)?(-5'sd12):(4'sd2)))));
  localparam [5:0] p2 = ((3'sd0)>(2'sd0));
  localparam signed [3:0] p3 = (~&{(^((-2'sd1)!==(2'd3))),((!(5'd22))===(~|(-5'sd1))),({(3'd6),(-5'sd8)}>={(3'd5),(4'd14)})});
  localparam signed [4:0] p4 = ((3'd4)<=(-2'sd0));
  localparam signed [5:0] p5 = ((((4'sd5)>=((-4'sd1)!=(-5'sd2)))|((4'd13)?(2'd2):(5'd5)))<=({1{((2'd2)?(3'd5):(5'd30))}}?((-3'sd2)?(2'd1):(3'd1)):((4'd9)?(2'sd1):(3'd4))));
  localparam [3:0] p6 = {4{{3{(4'd4)}}}};
  localparam [4:0] p7 = (-{{((6'd2 * (5'd26))!=(-4'sd5)),((~|(3'd7))^~(4'd2 * (2'd2)))}});
  localparam [5:0] p8 = ((5'd30)>=(-5'sd2));
  localparam signed [3:0] p9 = (~|{1{(&{2{{2{(^(3'd5))}}}})}});
  localparam signed [4:0] p10 = ((-4'sd0)?(4'd14):(2'd2));
  localparam signed [5:0] p11 = (~^{1{(^(~&(|({4{(2'd1)}}<((+(4'd1))|((4'd4)^~(2'd0)))))))}});
  localparam [3:0] p12 = {(2'd2),(5'd15)};
  localparam [4:0] p13 = ((((-2'sd1)?(5'sd8):(3'd1))?((2'd3)<(2'd1)):((3'd2)?(5'd25):(3'd3)))<<<{{3{(-5'sd7)}},((-2'sd0)-(-3'sd2)),(3'd3)});
  localparam [5:0] p14 = (((2'd3)?(4'd8):(3'sd1))?((3'd6)-(4'd5)):(~^(2'd3)));
  localparam signed [3:0] p15 = {((~(3'd7))^~(|(-2'sd0)))};
  localparam signed [4:0] p16 = (((3'sd0)^(4'd1))*((5'd22)===(4'd4)));
  localparam signed [5:0] p17 = {((5'd1)+(3'd0)),{(2'd2),(-3'sd2)},{(4'sd2),(4'd8)}};

  assign y0 = (($signed(($signed({4{$unsigned($signed(a3))}})))));
  assign y1 = (~^$unsigned($unsigned((|$signed((+$signed((^(~|$unsigned(((|$unsigned($unsigned((|(~&$signed(b3)))))))))))))))));
  assign y2 = ((a1^~b0)===(&(^a2)));
  assign y3 = (-5'sd6);
  assign y4 = ((5'd24)?((p3?p14:a3)==(p2>p16)):((p0?p4:p11)^(4'd15)));
  assign y5 = {(^(2'd1))};
  assign y6 = {4{(5'd8)}};
  assign y7 = {{3{p13}},{3{p13}},{(p11?p10:p15)}};
  assign y8 = {((p15?p12:p8)?($signed((p6?p15:p1))):{p16,p16,p15})};
  assign y9 = (-(^((4'd2 * {p2})+$signed(((|p13))))));
  assign y10 = (((p6||a1)>(p0<b1))^~((a2==a3)>>>(5'd20)));
  assign y11 = {1{((&p0)?(&p16):$signed(p7))}};
  assign y12 = (p4<<<p4);
  assign y13 = (&(!{(p15>>p4)}));
  assign y14 = {4{p9}};
  assign y15 = ((-((^(4'd2 * a0))>>>(~&(b0?b2:a5))))?($signed(((a5?a2:b4)?(-4'sd1):(a0||b1)))):{{a5,a4},(5'd2 * a1),{a2,a1,a0}});
  assign y16 = (5'd2 * (~^(+p1)));
  assign y17 = {(a5?b4:a4),{a5},(2'd3)};
endmodule
