module expression_00550(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((3'd6)?(5'sd6):(5'd10))?{(4'd14)}:((2'd1)?(5'sd12):(2'd0)));
  localparam [4:0] p1 = ((((2'd0)>(-2'sd0))>>((2'sd1)<<(3'sd2)))?(((3'd3)?(4'd4):(-5'sd15))&&{(5'sd14),(5'sd3),(4'd7)}):{(4'sd7),(4'sd6),(2'd3)});
  localparam [5:0] p2 = ((~^(2'd1))<<<(~(2'd3)));
  localparam signed [3:0] p3 = ({4{((-3'sd0)>(3'sd3))}}>((~((-4'sd7)&&(3'sd0)))!==((4'd13)^(4'sd6))));
  localparam signed [4:0] p4 = {3{((2'd0)>=(-5'sd11))}};
  localparam signed [5:0] p5 = ((-4'sd1)&(((2'd2)>>(3'sd3))>=((-2'sd0)===(4'd14))));
  localparam [3:0] p6 = ((((3'd0)?(5'd9):(3'd2))%(-2'sd0))-(4'sd3));
  localparam [4:0] p7 = {1{{1{{(((3'sd0)^(5'sd2))!={4{(5'd8)}}),(((5'd30)>>(2'd0))<<<{2{(3'd2)}})}}}}};
  localparam [5:0] p8 = (5'd2 * (-(^(3'd7))));
  localparam signed [3:0] p9 = ({3{(-3'sd3)}}<<{3{(2'd1)}});
  localparam signed [4:0] p10 = (((4'd2)<<<(4'sd7))>>{1{{4{(4'd3)}}}});
  localparam signed [5:0] p11 = ((~|((-4'sd6)>>(3'sd3)))!=={1{{1{(3'd1)}}}});
  localparam [3:0] p12 = ((~&(|(~|((2'd2)||(2'd3)))))<<<(~^((~|(5'd14))+((2'sd1)!=(-5'sd0)))));
  localparam [4:0] p13 = {{({2{(5'd8)}}?(~^(3'd3)):(~(-5'sd3)))},{{(-5'sd3),(2'd2),(5'd14)},(~&((5'sd13)?(5'sd4):(5'd19)))}};
  localparam [5:0] p14 = (~^(2'd3));
  localparam signed [3:0] p15 = (~|((!(2'd0))^~(|(5'sd2))));
  localparam signed [4:0] p16 = ((((-4'sd3)%(5'd7))||((5'd20)&(5'd27)))|(((-5'sd3)>>>(5'd22))+((5'd20)&&(4'd10))));
  localparam signed [5:0] p17 = {((+(4'd4))^(+(3'd7))),({(3'd7),(3'd3),(-5'sd8)}!=={2{(5'd11)}}),(!{3{(2'd0)}})};

  assign y0 = ((b3<<p11)*(b5==p5));
  assign y1 = (&(&(($signed((p17>=p6))>>>(p9>>p14))&&(~|((!(b3-a1))===((a1^~b4)))))));
  assign y2 = (a5!=p14);
  assign y3 = $unsigned($signed({1{a4}}));
  assign y4 = (|((^(b5>>b4))?{b1,b3}:(~{a0,a3,a5})));
  assign y5 = ($signed({3{p7}})-(2'd2));
  assign y6 = {2{(~^(+((b5&&a4)?(p6>a5):(a3>>>b5))))}};
  assign y7 = $unsigned($unsigned((~{1{(+b4)}})));
  assign y8 = {4{(b1|p13)}};
  assign y9 = {((b1!=p12)<(b3!==b2)),{(p11>p14),{3{p12}},(p1!=p5)},((p5+p6)&&{4{p2}})};
  assign y10 = (&((a1<=b0)!==(b4^b0)));
  assign y11 = {2{{{1{(p16?p9:p6)}}}}};
  assign y12 = (~^(|(+(~&(|(~|p5))))));
  assign y13 = (-(~((a1?b0:b2)?(-a2):(p11?b2:p13))));
  assign y14 = (!(+((a2!=b0)<<<(b0==b5))));
  assign y15 = ($unsigned($signed((3'sd0)))?$unsigned({2{(-5'sd14)}}):((4'd13)?{3{a1}}:(|p9)));
  assign y16 = $signed(((($unsigned(b1)=={1{a0}})<((p8^~p16)<<<(b0!==a1)))!={4{(~|(b0<p9))}}));
  assign y17 = {4{p1}};
endmodule
