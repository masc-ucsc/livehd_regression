module expression_00640(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd1);
  localparam [4:0] p1 = ({(2'd1),(3'sd0),(3'd2)}&((2'd3)>(5'd12)));
  localparam [5:0] p2 = (((~|(-4'sd0))<=((4'sd4)>>(5'd10)))?(+(-3'sd2)):(((-5'sd9)&&(2'sd0))+{3{(5'd6)}}));
  localparam signed [3:0] p3 = ((5'd7)^{4{(5'd17)}});
  localparam signed [4:0] p4 = (+((-4'sd2)*(-4'sd4)));
  localparam signed [5:0] p5 = ((4'd0)%(-4'sd3));
  localparam [3:0] p6 = (-4'sd7);
  localparam [4:0] p7 = (~|(3'd5));
  localparam [5:0] p8 = ((5'd21)>((3'sd3)!=(!(-2'sd1))));
  localparam signed [3:0] p9 = {2{(~((5'd9)||(4'd6)))}};
  localparam signed [4:0] p10 = {(2'd0),(-2'sd1),(-5'sd7)};
  localparam signed [5:0] p11 = ((-2'sd1)==(~|(~&(5'sd10))));
  localparam [3:0] p12 = ((((2'sd1)+(5'd15))!==((5'd30)&(2'd0)))==(((3'sd2)>>>(5'd15))+((5'd14)^~(4'sd2))));
  localparam [4:0] p13 = ({3{(3'sd2)}}>=(4'd9));
  localparam [5:0] p14 = ((((5'sd6)!=(-3'sd2))+((-3'sd3)?(2'sd1):(3'd3)))-({(3'sd2),(5'sd12),(3'sd0)}!=((3'sd3)?(4'sd7):(3'sd2))));
  localparam signed [3:0] p15 = (5'd2 * ((5'd19)<(3'd4)));
  localparam signed [4:0] p16 = (&(-2'sd0));
  localparam signed [5:0] p17 = ((5'd3)>>>(-2'sd0));

  assign y0 = (((b5>>>p15)?$signed(a3):(p16))&$signed((~^((b4?b0:p9)<{p15}))));
  assign y1 = ($unsigned((4'sd6))+(b2>>b0));
  assign y2 = ((((-p2)>=(a5!==a1))>((|b3)>(|a3)))>>(^{3{{2{p16}}}}));
  assign y3 = {1{(-5'sd9)}};
  assign y4 = {p6,p14};
  assign y5 = (3'd1);
  assign y6 = (((a0?p3:p10)?(p3?p13:a4):(b0<p15))^(+((~|(~|p15))%p13)));
  assign y7 = ({b2,p3}^~(p17?p10:p4));
  assign y8 = (2'd0);
  assign y9 = (2'd1);
  assign y10 = (~&(!(^{{4{b3}},(b3?a0:b3)})));
  assign y11 = (2'sd1);
  assign y12 = (-(p0?b1:b2));
  assign y13 = ($unsigned($signed(({(b2),(a4?a2:a4)}|((a5|a1)!=(a5?a5:b0)))))===(({a4,a5}^~(b3))<<<((a4>>>a3)||(a0<<b3))));
  assign y14 = (3'sd3);
  assign y15 = {{({p2,p13}!=(p17?a5:p13))},($signed(b0)?(a0<<<p2):(p0-p6)),((b3?b3:b5)===$unsigned((b4^a2)))};
  assign y16 = (a5?p9:b2);
  assign y17 = (-5'sd11);
endmodule
