module expression_00188(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd1)/(-3'sd1))<((-2'sd1)?(-2'sd1):(-2'sd0)));
  localparam [4:0] p1 = (&{4{{2{(3'd1)}}}});
  localparam [5:0] p2 = (|{((4'd9)&(5'd21))});
  localparam signed [3:0] p3 = (({((2'd2)<<(3'd3))}>>>(6'd2 * (3'd2)))<<<(3'sd3));
  localparam signed [4:0] p4 = ((-(3'sd0))^((4'd5)<<(3'd4)));
  localparam signed [5:0] p5 = {1{{4{(-5'sd2)}}}};
  localparam [3:0] p6 = (5'd0);
  localparam [4:0] p7 = {(((5'd5)?(2'd2):(5'sd13))+{4{(-3'sd1)}}),(|(-5'sd2))};
  localparam [5:0] p8 = {((-5'sd3)?(3'sd2):(4'd0)),{{(2'd1)},{(4'd11),(2'd0)}},((-3'sd3)?(5'sd7):(5'd6))};
  localparam signed [3:0] p9 = (~{{((|(3'sd0))?(~^(2'sd0)):{(3'd2),(3'sd3)}),{{(-5'sd15),(3'sd2),(-3'sd2)},{1{(3'sd2)}}}}});
  localparam signed [4:0] p10 = {(({(3'sd0),(-4'sd2)}^((4'd4)>>(4'd15)))>>>{((-4'sd6)!==(-2'sd0)),((5'sd3)>(-2'sd1)),(+(5'd23))})};
  localparam signed [5:0] p11 = {3{(4'd0)}};
  localparam [3:0] p12 = (~|(2'd2));
  localparam [4:0] p13 = (2'sd0);
  localparam [5:0] p14 = {(4'd1),{(4'd10),(3'sd3),(2'sd1)},((-5'sd7)?(-2'sd1):(5'sd15))};
  localparam signed [3:0] p15 = (3'sd1);
  localparam signed [4:0] p16 = {{(-5'sd14),(3'd2)}};
  localparam signed [5:0] p17 = {1{(^(~(!(-(^{3{(!(~^(-4'sd0)))}})))))}};

  assign y0 = {2{{2{p0}}}};
  assign y1 = (6'd2 * (a2+b2));
  assign y2 = (|(!((p6-p3)%p17)));
  assign y3 = (p3?p9:p9);
  assign y4 = {({3{a3}}!=(a5!=a4)),((-2'sd0)==(a1||a2)),((a4<<a1)||{(-3'sd2)})};
  assign y5 = (~|{1{p15}});
  assign y6 = $signed(({(a4&&a0)}<=(a3!==b0)));
  assign y7 = {3{({2{b3}}!==$signed({2{b3}}))}};
  assign y8 = (((p4%p17)/a3)==(4'd2 * (p2>>>p2)));
  assign y9 = (((!(&(a4+p2)))&(5'd2 * (a1==a1))));
  assign y10 = {2{p14}};
  assign y11 = (((p6))/a3);
  assign y12 = ((+$unsigned(p8))?(a0?a4:b1):(&{b3,a3,p7}));
  assign y13 = (((!p10)?(p2?b0:p7):(~|a4))?((p3?p4:p5)?(~&a1):(p0?p2:p10)):((p15?b4:p13)?(p9?p1:p8):(p16?p12:p1)));
  assign y14 = (({3{b1}}||{1{a4}})>>>$unsigned((~(a0?b1:b4))));
  assign y15 = (a3!==b3);
  assign y16 = (({b3,b4,b1}?{b5,a3,p17}:{a0})?({p3,a1,a0}?(b2>b1):{a5,a1,a4}):((a0?p11:p14)<<<(b1?a3:b5)));
  assign y17 = {(~(5'd22))};
endmodule
