module expression_00938(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd27);
  localparam [4:0] p1 = (5'd12);
  localparam [5:0] p2 = (~&(-5'sd12));
  localparam signed [3:0] p3 = ((&((5'd23)?(4'd13):(4'd12)))|(((-3'sd1)|(-2'sd1))>>((5'd26)?(3'd5):(2'sd0))));
  localparam signed [4:0] p4 = ({1{(~({1{((2'd2)<=(5'sd2))}}!==((2'sd1)^~(4'd0))))}}-((-((4'sd2)<(4'd6)))==((^(3'd0))==={4{(4'sd7)}})));
  localparam signed [5:0] p5 = ((((4'd12)?(3'd6):(5'd12))?((-3'sd1)+(4'd10)):((5'd19)!==(3'd0)))^(((3'd6)===(3'sd2))==((5'd16)||(4'd14))));
  localparam [3:0] p6 = ({3{(3'sd0)}}!==(-5'sd10));
  localparam [4:0] p7 = (+(^(4'sd0)));
  localparam [5:0] p8 = (3'd3);
  localparam signed [3:0] p9 = (!(-5'sd6));
  localparam signed [4:0] p10 = {(((2'd0)||(3'd0))+(~^(3'd6)))};
  localparam signed [5:0] p11 = (3'd7);
  localparam [3:0] p12 = {2{(((4'd6)==(-5'sd14))!==((2'd1)&&(3'sd3)))}};
  localparam [4:0] p13 = (-{2{(&(2'sd0))}});
  localparam [5:0] p14 = (4'd12);
  localparam signed [3:0] p15 = (-3'sd1);
  localparam signed [4:0] p16 = {1{(5'd2 * {(2'd0),(3'd1),(4'd12)})}};
  localparam signed [5:0] p17 = (((5'd7)?(3'sd3):(5'd8))>>((5'd13)?(3'd5):(5'd17)));

  assign y0 = ($signed((3'd2))!=(^(3'd5)));
  assign y1 = ({$unsigned({p11,b5,a5})});
  assign y2 = {2{{(p11?b3:p10),(p9>a4),{4{p15}}}}};
  assign y3 = ((+(!(!(+(a4^p16)))))&({2{b4}}^~{3{p16}}));
  assign y4 = ((b2?a3:a3)?(|(p12<<p4)):(b2&&a0));
  assign y5 = (&(&b4));
  assign y6 = (+((~^(p12<=p4))<<(3'sd0)));
  assign y7 = {{3{(b4>a1)}},{4{(b2&b0)}}};
  assign y8 = ({2{(a4||b4)}}>>>({b1}>(p0)));
  assign y9 = {4{(a1?p13:p11)}};
  assign y10 = (&((((p3?p1:p4)?(p11?p11:p11):(p13?p8:p8)))?($signed(p10)?(p14):(p2?p12:p7)):(-((|p7)?(p10):(p8?p4:p4)))));
  assign y11 = ({(p7!=p2),{p4,p1,p4},{p12,b1}}+({a2,a4}!==(b1^~a0)));
  assign y12 = (4'd14);
  assign y13 = $unsigned($unsigned($signed(((~&(({2{{2{b5}}}})))))));
  assign y14 = ((((a2!==b4)||{b3,a5,a5})<=((b3>>b3)===(a0<<a3)))!==$signed((4'd13)));
  assign y15 = ({p5,b4,a4}?{p0,p11}:(p8+p3));
  assign y16 = (|((~p2)?(&a5):(~|b0)));
  assign y17 = ((p9^~p7)?(p6?b1:p13):(b3?b3:p5));
endmodule
