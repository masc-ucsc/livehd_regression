module expression_00985(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-4'sd5)|(5'd2))<<((-3'sd3)^(5'sd7)));
  localparam [4:0] p1 = (6'd2 * ((3'd5)>=(2'd3)));
  localparam [5:0] p2 = (~&(!((~((4'sd0)^~(2'd0)))==(~|(4'd2 * (2'd1))))));
  localparam signed [3:0] p3 = ((4'd11)?(^(~&((3'sd3)?(3'sd1):(-2'sd1)))):(2'd2));
  localparam signed [4:0] p4 = {(2'sd1),(4'd6)};
  localparam signed [5:0] p5 = {(((-5'sd9)||(-3'sd0))^(&(-(2'sd0)))),(~&(^(((5'd0)>(3'd2))>(~|(-5'sd14)))))};
  localparam [3:0] p6 = (&(2'd2));
  localparam [4:0] p7 = ((-2'sd1)!=(&(((3'd7)*(5'd8))!=((-4'sd0)-(3'd3)))));
  localparam [5:0] p8 = {2{{2{(3'd6)}}}};
  localparam signed [3:0] p9 = (2'sd1);
  localparam signed [4:0] p10 = (((-2'sd1)?(3'd1):(5'sd1))/(2'd1));
  localparam signed [5:0] p11 = ((-((3'd2)?(3'd5):(4'sd2)))&&((4'd6)!=(-2'sd1)));
  localparam [3:0] p12 = {2{(4'd6)}};
  localparam [4:0] p13 = {(((-2'sd1)?(2'sd0):(-3'sd3))?((5'd8)?(2'd2):(-4'sd0)):{((2'sd0)?(-2'sd0):(4'd14))})};
  localparam [5:0] p14 = (+(6'd2 * ((5'd31)?(5'd0):(5'd17))));
  localparam signed [3:0] p15 = {(3'd0),(5'sd2),(2'd2)};
  localparam signed [4:0] p16 = {1{(5'd2 * {3{(3'd2)}})}};
  localparam signed [5:0] p17 = (({2{(3'd0)}}&&(+(2'sd1)))>>{4{(3'd0)}});

  assign y0 = $unsigned((~($signed(((-4'sd3))))));
  assign y1 = (~|(~&{(-3'sd3),(|($unsigned((4'd0)))),(+(4'd15))}));
  assign y2 = {((2'd2)&&(p14>>>b1)),{1{(3'd1)}},(-2'sd1)};
  assign y3 = ((a5)?(&p7):(~|b0));
  assign y4 = (p12<p16);
  assign y5 = (~{{b5},(4'd7),(4'd4)});
  assign y6 = {3{{a2,p4}}};
  assign y7 = $unsigned((~&{3{$unsigned((p15-p16))}}));
  assign y8 = ({4{p3}}?((a1?b3:a1)===(b4?b3:a0)):({1{b1}}!==(b2?a4:a2)));
  assign y9 = (!((5'sd14)|(3'sd0)));
  assign y10 = {{p15,a3,p10},(!b4),{a1,b4,b5}};
  assign y11 = (-3'sd1);
  assign y12 = {(3'd1),(5'sd3)};
  assign y13 = {2{((2'd0))}};
  assign y14 = (+(~(~|((~&(~^(-p4)))&&(+(p6>>>p11))))));
  assign y15 = (&a0);
  assign y16 = (5'd15);
  assign y17 = (({4{a5}}==(b2!==b2))||{3{b1}});
endmodule
