module expression_00085(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((4'd11)?(5'd21):(5'sd6)),((3'd7)?(-3'sd3):(5'sd3)),((2'sd1)?(4'd15):(4'sd2))};
  localparam [4:0] p1 = {2{{(5'd2 * ((5'd16)+(4'd5)))}}};
  localparam [5:0] p2 = (-4'sd7);
  localparam signed [3:0] p3 = (((2'd3)?(4'sd7):(-2'sd0))?((5'd25)?(2'd3):(-2'sd1)):{4{(4'sd7)}});
  localparam signed [4:0] p4 = ({(-5'sd11)}>=((3'd7)?(4'd13):(4'd10)));
  localparam signed [5:0] p5 = (^(~^({(4'd2 * (5'd3))}>>{{(5'd21),(-4'sd4),(-5'sd4)}})));
  localparam [3:0] p6 = (6'd2 * (5'd9));
  localparam [4:0] p7 = (-5'sd13);
  localparam [5:0] p8 = ((((2'sd1)?(3'sd1):(2'd0))?((2'd0)?(4'sd6):(2'd0)):((5'sd10)?(4'sd1):(5'd14)))!=(((5'd4)!==(3'd2))^((5'd25)-(2'sd0))));
  localparam signed [3:0] p9 = (+((5'd9)&(|(-3'sd2))));
  localparam signed [4:0] p10 = ((3'sd1)^(({2{(5'd5)}}-(2'd0))!=(|(-((-2'sd1)&(3'sd1))))));
  localparam signed [5:0] p11 = {(-3'sd3),(3'd6)};
  localparam [3:0] p12 = (4'sd6);
  localparam [4:0] p13 = ((4'sd4)<<{2{{4{(-4'sd7)}}}});
  localparam [5:0] p14 = {1{(~^{1{(((-5'sd3)||(2'sd1))^~(&(-3'sd2)))}})}};
  localparam signed [3:0] p15 = ((((-4'sd7)>>(3'd0))&&((-2'sd1)/(5'd0)))>=(((-4'sd5)!==(5'd19))-((4'sd2)==(4'sd7))));
  localparam signed [4:0] p16 = ({4{(3'd2)}}?{4{(2'sd0)}}:(2'd0));
  localparam signed [5:0] p17 = ((5'd30)!=(3'd4));

  assign y0 = {b4,p7,p4};
  assign y1 = (5'sd1);
  assign y2 = (~|{4{(~^{1{(b2<<a5)}})}});
  assign y3 = $unsigned({((+(5'd3))+((a5&&a3)?{b2,a0}:(p17^~b5)))});
  assign y4 = (~^(+({(p3),{p0,p4},{4{b0}}}?((a2?p4:p17)?(a5?p11:p8):(b3)):(^(~{4{b4}})))));
  assign y5 = (((a3?a5:b1)>(b2<=a1))?(2'sd1):((p3+p15)?(a3?b1:b2):(p0-p7)));
  assign y6 = (&(!((b0!==a1)*(~&b3))));
  assign y7 = (~&((+((3'sd3)==(a1?p1:p9)))?(4'sd2):((p13<p17)^(+a5))));
  assign y8 = ((({2{a1}}&(b4?a5:a1))>{2{(5'sd1)}})<=(^(2'd3)));
  assign y9 = {4{(!(|{3{p15}}))}};
  assign y10 = ((({p15}<<<(-p16))|((~&b2)==={b1}))^{((b4<b1)^~(a3+b3))});
  assign y11 = ({1{(b1<a5)}}<<<{3{a4}});
  assign y12 = ((&({(a4==b0)}))||({a2,b4}!==(b0)));
  assign y13 = ($unsigned({3{{a5,p14}}})?{(p7),(b1),(p0?a2:b5)}:{$signed(b5),{2{b2}},$signed(b3)});
  assign y14 = ({4{$unsigned((~|{2{b1}}))}});
  assign y15 = ($unsigned(((p0-p11)?{3{b5}}:(a3?p6:p0)))>=(($unsigned(a4)>>>(a5?p4:b5))-((p17+a2)>>>(a5?p13:b5))));
  assign y16 = {1{((&(+b2)))}};
  assign y17 = (!(^(+((&p3)+(+p5)))));
endmodule
