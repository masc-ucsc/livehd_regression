module expression_00402(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(^{(~|(3'd6)),{(3'd6)},{(-4'sd7),(-5'sd6),(4'd4)}}),{(-{(-2'sd1)}),(&(-(3'd7)))}}};
  localparam [4:0] p1 = ({(((5'd29)||(3'sd1))<{(4'd5),(5'sd4),(3'd4)})}>={(((5'd5)<(3'd2))+{{(-2'sd1),(-4'sd5)}})});
  localparam [5:0] p2 = ((5'd2)===(5'd22));
  localparam signed [3:0] p3 = {3{(4'sd5)}};
  localparam signed [4:0] p4 = (~^(~|({1{{((2'sd1)===(-4'sd6)),((5'd22)?(2'sd0):(3'sd0))}}}>>(~^({(4'sd4),(-3'sd1),(4'd8)}?{4{(4'd8)}}:(-(3'd4)))))));
  localparam signed [5:0] p5 = (((5'sd14)?(-5'sd15):(-4'sd7))?({4{(2'd0)}}||{1{(-3'sd0)}}):((3'd6)?(3'd2):(4'sd3)));
  localparam [3:0] p6 = {4{{3{(-5'sd9)}}}};
  localparam [4:0] p7 = (!((3'sd2)===(4'd0)));
  localparam [5:0] p8 = (~|(&{4{(3'd1)}}));
  localparam signed [3:0] p9 = {4{(5'sd15)}};
  localparam signed [4:0] p10 = ((-5'sd1)?(((-4'sd2)?(-4'sd1):(2'd1))+{3{(3'd7)}}):(-(4'd5)));
  localparam signed [5:0] p11 = ((~&(~&(-{3{(3'sd2)}})))?(!{2{{1{(5'd0)}}}}):(~&((-3'sd3)?(-3'sd0):(3'sd2))));
  localparam [3:0] p12 = {2{({4{(-5'sd12)}}?((5'sd8)+(5'd12)):(&(4'd14)))}};
  localparam [4:0] p13 = (4'sd1);
  localparam [5:0] p14 = (|{3{(~&(&(4'sd7)))}});
  localparam signed [3:0] p15 = (((~|(5'd3))+((-4'sd7)/(5'sd8)))-(((3'd1)!==(4'sd6))*((3'd7)%(4'd12))));
  localparam signed [4:0] p16 = (~((-(&(!(!(3'd5)))))&&((2'd0)||(-3'sd0))));
  localparam signed [5:0] p17 = (((((4'd1)>>(3'sd1))>((5'sd11)||(-5'sd3)))==(6'd2 * ((4'd8)<<<(3'd2))))^~(5'd2 * ((5'd31)==(4'd11))));

  assign y0 = {(&p13),(~p15)};
  assign y1 = $unsigned($unsigned($unsigned(({b5,b3}!==(b0===b3)))));
  assign y2 = {3{{{p2},{2{b0}}}}};
  assign y3 = (~($unsigned(p5)<<{a5}));
  assign y4 = (~|(((b1!=b0)<=(a5?b5:a0))?{3{b4}}:(+{1{{a4,b5}}})));
  assign y5 = (~((3'sd1)!==(5'd4)));
  assign y6 = $signed((((b3?b2:b0)^(b4?a0:b0))<<($signed((b5?p4:a1))*$signed((b0?a0:b3)))));
  assign y7 = (b1<b2);
  assign y8 = ((-5'sd14));
  assign y9 = $signed((((4'd0))>>((a4?b5:a2)?(b0>>a2):(-5'sd0))));
  assign y10 = {{4{(-3'sd0)}}};
  assign y11 = (3'd6);
  assign y12 = {3{({3{p11}}>=(p12&p16))}};
  assign y13 = (((b4==b0)>=(a0))===(&$signed((~&(b4===a2)))));
  assign y14 = (-(((|a3)<(^p9))-(&(2'd1))));
  assign y15 = (p14?b4:a5);
  assign y16 = {{(a3?p9:b3),(p10?a2:a1),(p16?p1:p14)}};
  assign y17 = (-2'sd1);
endmodule
