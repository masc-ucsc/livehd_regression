module expression_00469(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+((4'sd4)?(|((4'd13)==(3'sd2))):(|(+(2'd3)))));
  localparam [4:0] p1 = {{(-2'sd0)},{(4'd0)}};
  localparam [5:0] p2 = (~|(2'sd1));
  localparam signed [3:0] p3 = {(5'd0),(&(~&((5'd29)<<(4'd11)))),((^(2'd0))<<{(2'sd1),(2'd1)})};
  localparam signed [4:0] p4 = (5'd22);
  localparam signed [5:0] p5 = (+{({(2'sd1),(3'd2),(-2'sd0)}<<<{(3'sd2),(3'sd0)}),(~|{((4'd0)-(4'sd4)),((4'd13)|(5'd30))}),(+((&(4'sd1))>>>((2'd0)===(3'd0))))});
  localparam [3:0] p6 = {3{{1{(3'd0)}}}};
  localparam [4:0] p7 = (~|(~&({4{(4'sd7)}}^~(^(2'sd1)))));
  localparam [5:0] p8 = ((^{3{(5'd5)}})===(4'd12));
  localparam signed [3:0] p9 = (((4'd14)!==(2'd0))<<(|((2'd2)%(-2'sd0))));
  localparam signed [4:0] p10 = ((((-3'sd1)>=(2'd3))||((3'sd2)>>>(-3'sd3)))>(+((!((2'd1)>(4'd5)))>>>((4'd0)<<<(2'd1)))));
  localparam signed [5:0] p11 = ((((4'd4)<(2'sd0))?((-2'sd1)?(4'sd4):(-5'sd9)):((4'd11)<<<(3'd6)))?(~|(-((4'd2)===(2'd2)))):(-2'sd0));
  localparam [3:0] p12 = ((((4'sd6)<=(2'd1))||{2{(2'd3)}})?(((3'd5)|(3'd5))<=((5'sd10)!=(2'd0))):((2'sd1)?(-3'sd0):(5'd7)));
  localparam [4:0] p13 = ((4'd3)?(2'd1):(3'sd0));
  localparam [5:0] p14 = (({(-4'sd5),(5'sd7),(-5'sd7)}>((3'd4)>>(3'd2)))>>>((~^(~(2'sd0)))>>(&((5'sd3)>(4'd14)))));
  localparam signed [3:0] p15 = ((^{4{(4'd15)}})>((~|((2'd2)&&(2'd2)))=={1{(2'd3)}}));
  localparam signed [4:0] p16 = (!(-3'sd0));
  localparam signed [5:0] p17 = ({{3{(4'sd6)}},((3'd0)<(5'd5)),(~|(2'sd1))}<<<(~|(+(((2'sd1)<<<(-3'sd0))!==(+(3'd4))))));

  assign y0 = (&(&(^p1)));
  assign y1 = {4{{1{a1}}}};
  assign y2 = (p11?p10:p2);
  assign y3 = (2'd2);
  assign y4 = (-5'sd13);
  assign y5 = (^{3{((+p5)?(p17!=p14):(p12==p10))}});
  assign y6 = {((p13-p3)<(a4^~p0)),{(p16&b3),(b3?p6:p2),(p8?p9:p3)}};
  assign y7 = {(4'd2 * b2),{a5,b5}};
  assign y8 = (-4'sd0);
  assign y9 = (+{(~^{b5}),{a1,a4,a1}});
  assign y10 = {({4{(+p4)}}<<(-{1{{1{{1{{1{{2{a0}}}}}}}}}}))};
  assign y11 = (($unsigned(p14)<=(b2?p12:b5)));
  assign y12 = (5'sd14);
  assign y13 = {{{(~|(~|p11)),{a4,p1,b0}},(!{{b5},{a1}}),(-(|{{p17,p13},(|a3)}))}};
  assign y14 = ({((p17?p12:p8)?{3{b4}}:{2{p16}})}==((p13!=p10)?(p8?b0:p14):(a5==b5)));
  assign y15 = (a4|p12);
  assign y16 = ((~^(p3|p1))%p15);
  assign y17 = (-4'sd5);
endmodule
