module expression_00002(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (2'd1);
  localparam [4:0] p1 = {(3'd0),(3'd7)};
  localparam [5:0] p2 = (5'd10);
  localparam signed [3:0] p3 = {((4'd15)?(2'sd0):(4'sd3)),(((4'd15)^(5'd31))|((5'd27)?(3'd5):(2'd1))),((4'd5)?(4'd7):(5'd21))};
  localparam signed [4:0] p4 = (^((-5'sd0)<=(2'd2)));
  localparam signed [5:0] p5 = ((((5'sd15)|(4'd11))==((3'd0)?(3'd7):(-5'sd4)))&({4{(3'd2)}}=={1{((3'd5)?(4'd11):(4'd13))}}));
  localparam [3:0] p6 = (-(((~((-4'sd6)>(-3'sd1)))!==((3'd5)<<(5'sd0)))!=(5'd0)));
  localparam [4:0] p7 = {2{(!(~{3{(-5'sd9)}}))}};
  localparam [5:0] p8 = ((((-4'sd4)+(2'sd1))<((4'sd5)&(5'sd10)))<((4'd2 * (4'd13))&((-2'sd0)<<(5'd3))));
  localparam signed [3:0] p9 = {{(-3'sd1),(3'd1),(4'sd3)},{(2'd1),(-4'sd1),(5'sd15)}};
  localparam signed [4:0] p10 = {(~|((2'd3)?(4'd11):(4'd9))),(~^{1{((3'd1)?(3'd1):(5'd14))}})};
  localparam signed [5:0] p11 = ({3{(3'd4)}}?({2{(5'sd9)}}^~{(5'sd9),(4'd3),(-5'sd3)}):(((2'd1)>>(-4'sd0))-((5'd2)?(2'sd1):(3'd0))));
  localparam [3:0] p12 = ((((5'sd0)^~(4'sd6))!==((3'sd3)<<(-5'sd5)))?(-((5'd6)?(4'd15):(-5'sd8))):(5'd6));
  localparam [4:0] p13 = ((3'sd2)?(-5'sd5):(5'd1));
  localparam [5:0] p14 = (~^(!{{(-2'sd1),(-5'sd8)},(~|((4'd7)<(4'd3))),(!{(-4'sd6),(3'sd0),(4'sd0)})}));
  localparam signed [3:0] p15 = (((5'd11)&(-4'sd5))^((5'sd4)<<(2'd1)));
  localparam signed [4:0] p16 = {3{((2'd1)<(3'sd1))}};
  localparam signed [5:0] p17 = ({3{(2'd0)}}?((3'd0)?(-5'sd1):(2'sd1)):(((-3'sd0)===(3'sd0))-((3'd3)===(5'sd14))));

  assign y0 = ({((4'd15)===({4{b3}}>>>(a4==a1)))}!={3{(p9<=p14)}});
  assign y1 = ((6'd2 * p0)^(2'sd1));
  assign y2 = {2{(({3{b0}}!=(p6==p1))!={1{{1{(5'd30)}}}})}};
  assign y3 = ({4{b1}}?{4{a5}}:{1{{4{b2}}}});
  assign y4 = $unsigned((&(^$unsigned((+$signed($signed(a1)))))));
  assign y5 = (+(p6?p3:p14));
  assign y6 = (-(b3<b4));
  assign y7 = ((3'sd3)<<<((-2'sd0)));
  assign y8 = ((!(((b1-a5)&&(a1!==b0))===(|(b1&b1))))<<<((^(!(a0<<p12)))>=((a4^a5)!==(b5!==b5))));
  assign y9 = ((~$unsigned({(b3),(a5?a0:a5),{3{b4}}}))?{4{(a3?p8:a2)}}:$unsigned((~|{4{a1}})));
  assign y10 = (~|((~(~(-p10)))^(-(-(p4||a4)))));
  assign y11 = ({a5,b1,a1}==(5'd24));
  assign y12 = (((-4'sd4))^(((p2+b2)==(4'sd3))|((a0==b1)==(2'sd0))));
  assign y13 = ((b2<b0)==(p7>=p6));
  assign y14 = {((5'd2 * (-(+b2)))<<$signed({(b5>>p8),{p4,p16}}))};
  assign y15 = $signed((-(~({2{b2}}?$signed((b5-b1)):(p5>>>a0)))));
  assign y16 = $unsigned((~^(3'd2)));
  assign y17 = (~&(5'd14));
endmodule
