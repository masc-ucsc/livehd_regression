module expression_00740(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{{1{(5'd21)}},{(2'd3),(3'd0)}}}};
  localparam [4:0] p1 = (^(!(2'd0)));
  localparam [5:0] p2 = {((2'd2)<(3'd4)),((3'sd2)<<(2'sd0)),((5'd25)>(2'sd0))};
  localparam signed [3:0] p3 = (((2'd0)?(3'd7):(-5'sd5))?{{(-2'sd0),(2'd3)}}:((-5'sd10)?(3'd6):(3'd5)));
  localparam signed [4:0] p4 = (~((~^((-3'sd2)?(3'd2):(-3'sd3)))?((4'sd2)?(-3'sd3):(2'd2)):((5'd11)?(-3'sd3):(5'sd12))));
  localparam signed [5:0] p5 = ((4'd9)!==(5'd8));
  localparam [3:0] p6 = (((4'd6)<=(3'd5))?((-5'sd12)==(5'd26)):(4'd15));
  localparam [4:0] p7 = ((2'sd0)==(-2'sd1));
  localparam [5:0] p8 = (((2'd3)^~(3'd0))|((5'sd6)<=(-2'sd1)));
  localparam signed [3:0] p9 = (~(~&(^(5'd20))));
  localparam signed [4:0] p10 = {{{(4'd12),(2'd0)},{(2'd3),(5'sd8)},((4'sd6)-(5'd3))}};
  localparam signed [5:0] p11 = {((-5'sd3)|(2'sd1)),((-5'sd0)<=(4'sd7))};
  localparam [3:0] p12 = (-5'sd9);
  localparam [4:0] p13 = ((((-4'sd4)!==(3'sd0))===((5'd18)+(-4'sd4)))<<<(((5'd21)-(4'd10))|((5'd16)!=(4'd5))));
  localparam [5:0] p14 = {2{((4'sd3)^~{3{(-4'sd4)}})}};
  localparam signed [3:0] p15 = {(5'd23),(3'd5),(~&(4'sd1))};
  localparam signed [4:0] p16 = ({{(-3'sd1),(3'd2),(3'd7)},((4'd15)?(2'sd1):(5'd1)),(!(2'd3))}>>>(((4'sd4)?(3'd4):(2'd1))?{(3'sd2)}:{(-2'sd1),(2'd0)}));
  localparam signed [5:0] p17 = ((5'd21)?((2'd0)?(4'd12):(5'sd12)):((3'd6)?(5'sd0):(4'd4)));

  assign y0 = (3'd0);
  assign y1 = (+{{4{{a3,a0,b3}}},{{1{a2}},(2'd2),{1{b2}}}});
  assign y2 = $unsigned((((a5>=p9)&(~^p11))));
  assign y3 = ((^{2{{b1}}})?{{{2{{a1,p15,p9}}}}}:((p8?b4:p17)!=(&(a5===b1))));
  assign y4 = (({2{a4}}?(a4>>>p5):$signed(p4))?$unsigned(((p12?p14:p6)-(a4===b0))):((+{4{a4}})));
  assign y5 = ((p3?p14:a1)<=(4'd2 * p1));
  assign y6 = (((~|{2{p15}})=={4{p8}})<<<(~&((p11<<b4)<<{p15,a4})));
  assign y7 = ({(^p5),(~b3),(~&b2)}?(!{1{{{a1,b1}}}}):(^{(p6?a5:b2)}));
  assign y8 = (-5'sd8);
  assign y9 = (^a2);
  assign y10 = (|({1{((-$unsigned(((^(~|a0))?(^$unsigned(a2)):{3{b1}}))))}}));
  assign y11 = (2'd1);
  assign y12 = (((p11)>=(b1^a2))||$unsigned({3{a5}}));
  assign y13 = $signed({4{a4}});
  assign y14 = (5'd13);
  assign y15 = {b4,b5,p16};
  assign y16 = {2{{2{(b1?b2:a2)}}}};
  assign y17 = ((b5^~p10)*(~^(a1>a5)));
endmodule
