module expression_00209(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (+(3'sd3));
  localparam [4:0] p1 = (4'd2 * (^((4'd9)>(3'd4))));
  localparam [5:0] p2 = (((((-4'sd7)!==(5'd15))-((3'd5)&(2'd0)))!==(|(|((5'd12)===(3'd6)))))==(~(^((~((3'd2)-(4'd9)))^~((-5'sd12)|(3'd7))))));
  localparam signed [3:0] p3 = (~^(({(-3'sd0),(5'sd10)}!=((3'd6)|(3'd6)))-{((3'd2)<<<(5'sd0)),{(-2'sd0),(3'sd1),(-4'sd7)},(&(4'd14))}));
  localparam signed [4:0] p4 = (^(-5'sd1));
  localparam signed [5:0] p5 = (2'd1);
  localparam [3:0] p6 = (((4'sd6)+(5'd0))/(4'd9));
  localparam [4:0] p7 = {(-4'sd6),(3'd3)};
  localparam [5:0] p8 = (3'sd3);
  localparam signed [3:0] p9 = {3{(-2'sd0)}};
  localparam signed [4:0] p10 = ({(5'd22),(-4'sd1)}==((-5'sd2)<(3'd3)));
  localparam signed [5:0] p11 = (4'sd4);
  localparam [3:0] p12 = {(((2'sd0)-(4'sd6))&&{3{(5'sd2)}}),{2{{(5'd17),(-4'sd3)}}},{4{(3'd6)}}};
  localparam [4:0] p13 = (({(-4'sd4),(5'd18),(3'd0)}?((-4'sd1)-(5'd2)):{(4'sd1),(5'd7)})-(((5'd22)?(-4'sd5):(2'd1))?{(5'sd3),(3'sd1)}:((2'd1)==(5'sd9))));
  localparam [5:0] p14 = {(-2'sd0)};
  localparam signed [3:0] p15 = (!(-(&(~&((4'sd2)>>{1{(-2'sd1)}})))));
  localparam signed [4:0] p16 = {(5'd14),((!(-4'sd5))?((2'sd1)!==(-4'sd6)):(-5'sd12))};
  localparam signed [5:0] p17 = ((^({2{(2'd2)}}<={2{(4'd11)}}))|{4{((3'd2)?(4'd15):(4'sd0))}});

  assign y0 = {4{(~&(a0+b5))}};
  assign y1 = ((p3^~p10)<(5'd2 * p12));
  assign y2 = {(4'd2),{{b2},{p1,a2},(b5?p9:p1)},{(5'sd15)}};
  assign y3 = (~|(((!(b0<b0))<<(2'd3))>>(2'd0)));
  assign y4 = {({b2}?(2'd2):{1{p9}}),({3{b0}}?{a1,p14}:{a3,p9}),((2'sd1)?{a5,p2}:{4{b5}})};
  assign y5 = ({(a3-a1),(a0!=b4),(a1^a3)}&&(-3'sd1));
  assign y6 = ($signed(($unsigned((a1?b0:b3))))^$signed(((a1)>=$signed(a1))));
  assign y7 = ({2{p2}}!=(p2>>a3));
  assign y8 = (((~|((5'd22)))>>{4{p17}})>(5'd10));
  assign y9 = (+((4'd14)&&(2'd3)));
  assign y10 = (~|{2{((|(p0^a4))^~(^(p11?p5:p15)))}});
  assign y11 = (~|{3{(p5&a2)}});
  assign y12 = (((b5!=p11)?{4{p9}}:(p2^~p10))<<((~^p5)<{p12,p15}));
  assign y13 = (((3'd4)?(a4?a1:a0):(|p5))<=(!((b0!==a2)<<<(4'd15))));
  assign y14 = {3{(p4!=p9)}};
  assign y15 = ((~|((a0>b2)?(b0>=a3):(b2)))<((5'sd3)?(a0>>>b3):(a5!=a5)));
  assign y16 = (+{2{{2{b2}}}});
  assign y17 = (~^(!(((^p2)>>>(4'd3)))));
endmodule
