module expression_00436(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {4{(3'd7)}};
  localparam [4:0] p1 = ((~((5'd30)?(-5'sd4):(4'd11)))?(~|((4'd0)?(-5'sd5):(2'd3))):((~|(-4'sd4))*(-(-3'sd0))));
  localparam [5:0] p2 = (4'd6);
  localparam signed [3:0] p3 = ((!((~|((5'sd13)<<<(5'd14)))>(~&((4'd0)*(2'sd1)))))==(~&(~&(((2'sd0)||(3'sd2))<<<((2'sd0)!==(3'd2))))));
  localparam signed [4:0] p4 = {1{({3{(&(4'd3))}}>>>(~&{4{((2'sd0)>=(-5'sd11))}}))}};
  localparam signed [5:0] p5 = (4'd4);
  localparam [3:0] p6 = ({1{((5'd5)&&(4'sd1))}}^{3{(-3'sd2)}});
  localparam [4:0] p7 = (~&{2{(-3'sd1)}});
  localparam [5:0] p8 = ((((2'sd1)?(3'd5):(2'd0))^~((2'd3)?(3'd4):(2'sd0)))>={3{((5'd12)>=(-4'sd1))}});
  localparam signed [3:0] p9 = {3{((4'sd0)>(5'sd8))}};
  localparam signed [4:0] p10 = (((-2'sd0)==(4'd9))===((2'sd0)>>>(3'd0)));
  localparam signed [5:0] p11 = {((~^(5'sd1))?(|(3'sd3)):{3{(-4'sd6)}})};
  localparam [3:0] p12 = {2{(~|{4{((5'd22)^~(-3'sd3))}})}};
  localparam [4:0] p13 = {{1{(4'd4)}},{(4'sd6)}};
  localparam [5:0] p14 = {3{{1{(-3'sd3)}}}};
  localparam signed [3:0] p15 = ((~(((5'sd7)<(3'sd1))!=(~&(2'd1))))>>>{(-(4'sd1)),((-5'sd1)&&(5'sd1)),((2'd1)>>(3'sd1))});
  localparam signed [4:0] p16 = (+((~&(((4'sd2)?(2'd1):(5'sd12))^~((4'd3)?(4'sd1):(4'd14))))<=(~^({(2'd3)}?{(3'd6),(2'd1)}:(~^(3'd0))))));
  localparam signed [5:0] p17 = {2{(((4'd15)&&(3'd6))<=((-2'sd0)!==(-5'sd10)))}};

  assign y0 = (((b3!=a0)&{p0,a1,b3})^((p11?p6:p3)^~(a4&p17)));
  assign y1 = ((p6||b5)^(b2||a2));
  assign y2 = (((p10>p3)*(p12&p3))?((p0>>>p12)&(3'd1)):((p14<<p8)?(p5?p11:p9):(p16?p11:p17)));
  assign y3 = (((2'd2)%p7)==(^(4'd0)));
  assign y4 = (((b5>>p16)<(-2'sd1)));
  assign y5 = ($unsigned((($unsigned((p5?p8:b1))>{p13,p13})?({a4,b2}<<<{a1,p16,a3}):({(p4?p6:p17)}>=(p6?p8:p5)))));
  assign y6 = ((2'd3)==((|p0)?(+p0):(p12&&p9)));
  assign y7 = (b4-b4);
  assign y8 = {1{{1{((-4'sd6)>>>{(3'd1),{p1}})}}}};
  assign y9 = {(!{{a5},(a0===a5)}),{{p4,p0},$signed((b5<<<a0))},((!$signed(a3))>={{2{p2}}})};
  assign y10 = ({b1,p9,p12}||(p1&&a2));
  assign y11 = ((p0&p6)>>(p1-a1));
  assign y12 = (^{4{(~^p9)}});
  assign y13 = ((3'd1)===((2'd1)!==(a2?b1:a3)));
  assign y14 = (((b5===b5))?(a0+p2):$unsigned((p12)));
  assign y15 = ((-{4{(p3^~p5)}})<<{{a2,b2,a1},{3{a4}},{p8,p4}});
  assign y16 = (~^{(4'sd5),(-p3),(+p16)});
  assign y17 = (({(b4^a4)}!==((a5>>>b0)^~(5'd2 * a2)))&&{{(3'd3),{a2,a3,a4},(4'sd5)}});
endmodule
