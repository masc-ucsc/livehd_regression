module expression_00702(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((2'd0)|(4'sd2))+(!((-3'sd3)<<<(-3'sd0))))};
  localparam [4:0] p1 = ((3'd7)?(-2'sd0):(2'sd1));
  localparam [5:0] p2 = {2{(~^{((4'sd2)?(4'sd7):(5'd18)),((4'd11)?(-4'sd2):(3'd6)),{4{(-5'sd3)}}})}};
  localparam signed [3:0] p3 = (((3'sd3)>>(5'd18))<=((-5'sd13)!==(5'd17)));
  localparam signed [4:0] p4 = (5'sd13);
  localparam signed [5:0] p5 = (({3{(5'd25)}}==(6'd2 * (3'd3)))||{(~&(5'd22)),((3'sd0)>=(-4'sd4))});
  localparam [3:0] p6 = ((((-2'sd1)^(-3'sd2))<={(4'd15),(4'd11),(2'd2)})?(((-2'sd1)?(2'd0):(-2'sd0))?((-3'sd3)!==(-3'sd1)):((3'd5)?(-5'sd6):(4'sd4))):(((-2'sd0)&&(2'd1))>{(5'd0),(5'd14)}));
  localparam [4:0] p7 = (-(4'd14));
  localparam [5:0] p8 = (5'd14);
  localparam signed [3:0] p9 = ((~(+((&(5'sd14))|(^(3'd6)))))&&(+(~(((4'd2)<<<(5'd31))==((4'sd6)&&(2'd3))))));
  localparam signed [4:0] p10 = (4'd13);
  localparam signed [5:0] p11 = (3'd6);
  localparam [3:0] p12 = {4{{(5'sd3),(-3'sd3)}}};
  localparam [4:0] p13 = {(((3'd1)===(3'd5))&((5'd19)^(3'd6))),{(((3'd3)+(3'd2))<<{(3'd2),(4'd14)})}};
  localparam [5:0] p14 = {(5'd7),(3'sd2),(2'd0)};
  localparam signed [3:0] p15 = ((((5'sd4)^~(2'sd1))|((3'sd0)-(2'sd0)))^~{(^(-5'sd3)),(+(2'd3))});
  localparam signed [4:0] p16 = (&{(&(~^{4{(5'd2)}})),{{{(4'sd2)},{(3'd7),(5'sd9)},{(3'd4)}}}});
  localparam signed [5:0] p17 = ({((-5'sd13)>>(5'd17)),(|(3'd4)),(!(5'd8))}?(+((&(3'd5))!==((5'd19)|(-2'sd0)))):(((3'sd0)&&(2'd2))?(~&(3'sd1)):{(-2'sd0)}));

  assign y0 = {a1};
  assign y1 = (5'sd13);
  assign y2 = (~&(({2{p11}}>{3{b2}})&((-3'sd1)<<(-(a0!==b2)))));
  assign y3 = $unsigned(((p10<<p14)>=(a5<<<b4)));
  assign y4 = ((^((a1<<b1)===(b5*b0)))+((p14>>>b0)|(b3<=p16)));
  assign y5 = ({(~&{2{(p4!=a1)}})}<<<$signed(((-(|p6))+(a0!=p8))));
  assign y6 = (~((((~&p2)/p6)&&(-(b4!=p14)))>>>(((p10%p17)==(|p10))<<<((~b3)<(p16!=p8)))));
  assign y7 = {(+(5'd2 * (5'd15))),{(4'd2 * b2),(5'd17),(a3>>a5)}};
  assign y8 = {2{(5'd7)}};
  assign y9 = (({1{p17}}|(p5<<p2))=={1{{2{p6}}}});
  assign y10 = ($unsigned(((b2?a0:a5)?(~|(a2?b0:b3)):(&(|b0)))));
  assign y11 = {(a0?a3:p16),(-4'sd4),(b5^~b0)};
  assign y12 = ((a5|b5)?{p0,b4}:{p14,p3,b0});
  assign y13 = {3{((p17^p0)?(~^a1):{p17,p4,b0})}};
  assign y14 = ((!(p1>=p0))<=(3'd3));
  assign y15 = ((({(b2<b2)}<<$signed((a2&b0))))<<<{{((b4?a5:b0)>(b3)),(b5?p1:a4)}});
  assign y16 = (2'd3);
  assign y17 = (!(2'd2));
endmodule
