module expression_00858(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((&((5'd22)>=(2'd1)))*(|((3'd6)?(-4'sd3):(-3'sd0))));
  localparam [4:0] p1 = (-3'sd3);
  localparam [5:0] p2 = (&(3'sd1));
  localparam signed [3:0] p3 = {{{(-3'sd0)},(!(-2'sd0)),(-5'sd6)},({(-4'sd3),(-2'sd1)}?{(-5'sd5),(4'sd6)}:(3'd2)),{2{(~&(4'd9))}}};
  localparam signed [4:0] p4 = {(2'd1),(3'd2),((4'sd1)|(2'd0))};
  localparam signed [5:0] p5 = ({(((-2'sd1)<(-4'sd2))||(-2'sd1))}>=(3'd5));
  localparam [3:0] p6 = (|(~|(|(!(+(+(-2'sd0)))))));
  localparam [4:0] p7 = (~&((4'sd4)?(5'd11):(2'd1)));
  localparam [5:0] p8 = {{((2'd2)<<<(2'd3))},{((5'd27)<=(5'sd0))},((2'sd0)&(-2'sd0))};
  localparam signed [3:0] p9 = ((~^(+(4'd9)))^{4{(5'd9)}});
  localparam signed [4:0] p10 = {{{(~|{(~{(-5'sd8),(2'd1)}),(~^{(4'd13),(4'd6),(5'd9)})})}}};
  localparam signed [5:0] p11 = (|(5'd0));
  localparam [3:0] p12 = (4'd9);
  localparam [4:0] p13 = ((&(-(-(-3'sd1))))?((-5'sd13)?(3'd7):(-3'sd3)):(&{2{(3'sd2)}}));
  localparam [5:0] p14 = {4{((3'sd1)^~(-2'sd0))}};
  localparam signed [3:0] p15 = {((4'd4)!==(-3'sd2)),(^(5'sd12)),((2'd1)>=(-2'sd1))};
  localparam signed [4:0] p16 = {3{((-4'sd0)<<<(3'd6))}};
  localparam signed [5:0] p17 = {2{(((3'd6)>=(-5'sd4))>(&(2'sd0)))}};

  assign y0 = (3'sd1);
  assign y1 = ((^b5)<(b2<a1));
  assign y2 = (-((p5?p12:p8)>=(!a3)));
  assign y3 = ((|(~a1))<<(+(~^b5)));
  assign y4 = (4'd12);
  assign y5 = ((-3'sd2)>((a2/p17)?(p11<a4):(p9==p2)));
  assign y6 = {({((~(5'd2 * p12))?(p11?p16:p8):(|{p11,p13}))}+{(p10?p16:p14),((p3?p3:p8)<<<(!p1))})};
  assign y7 = $signed(((+(|(2'd2)))!=({$signed((-2'sd1))}&&($unsigned(b5)!=={a3,b1,a2}))));
  assign y8 = {2{(b5>>>a4)}};
  assign y9 = ((p13?p1:a5)?(5'sd10):{2{b1}});
  assign y10 = (((a4?a5:b1)===(|a1))?({1{p7}}|(p4-p2)):((p17>=p1)?(2'sd1):(p17|p3)));
  assign y11 = ((p14<=p5)-(b3!==b0));
  assign y12 = $unsigned((-((b2?b2:p11)==(a2^p14))));
  assign y13 = (4'd2 * {3{a2}});
  assign y14 = {3{(-2'sd0)}};
  assign y15 = ((~(p11+p5))?(!(a0===a5)):(p13<<<p13));
  assign y16 = {3{(5'sd8)}};
  assign y17 = (~(3'd7));
endmodule
