module expression_00043(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(5'd12)};
  localparam [4:0] p1 = ({({3{(2'sd0)}}&&((5'd18)<(-2'sd0)))}+(((3'd6)?(5'd10):(5'sd11))>>({(5'sd6),(2'sd0),(2'sd0)}-((5'd29)==(-3'sd1)))));
  localparam [5:0] p2 = (((2'sd0)/(5'sd11))*((-4'sd7)<<<(3'd7)));
  localparam signed [3:0] p3 = (+(-({(3'sd2)}>{(-4'sd4)})));
  localparam signed [4:0] p4 = (((4'sd5)&(5'd9))?((-3'sd0)&&(5'd30)):((3'd4)<<<(3'd7)));
  localparam signed [5:0] p5 = ({4{(2'd1)}}<<(((-2'sd1)>=(3'd0))&((5'sd8)^(5'd29))));
  localparam [3:0] p6 = ((-3'sd2)&(2'd3));
  localparam [4:0] p7 = (~^{{(^(|(2'd1))),(&(^(4'd15)))},((+{(4'd8),(2'sd0)})-((2'd2)?(-4'sd2):(-5'sd4)))});
  localparam [5:0] p8 = (({4{(-5'sd7)}}<<(~|(4'sd1)))<=(~&{3{(-3'sd1)}}));
  localparam signed [3:0] p9 = {((5'sd15)+(4'd7))};
  localparam signed [4:0] p10 = ({(-5'sd5),(-2'sd1),(4'd15)}>>{(3'sd1),(4'd10),(3'd3)});
  localparam signed [5:0] p11 = (((-4'sd1)>>(3'sd2))^~((-5'sd9)===(4'd11)));
  localparam [3:0] p12 = ((4'd13)>(2'd1));
  localparam [4:0] p13 = (~|{((2'd2)?(4'sd3):(4'd9)),(~(-{(4'sd1)})),(!{(-3'sd1),(-3'sd3)})});
  localparam [5:0] p14 = (((3'sd2)||(5'd26))>>{1{(&(-5'sd3))}});
  localparam signed [3:0] p15 = {{{(-2'sd0),(-2'sd1)},{(3'd4),(4'd3)},{(-2'sd1),(-5'sd5)}},{{(4'd3)},{(2'd3),(3'sd2)}},{{(4'd9)},{(3'sd0),(-5'sd8)},{(-4'sd2),(2'd3),(-5'sd7)}}};
  localparam signed [4:0] p16 = (^(+(2'sd1)));
  localparam signed [5:0] p17 = (~&(~&(((3'd5)>>>(-4'sd3))<<((3'd7)>>>(5'd30)))));

  assign y0 = (~^(p9?p9:p14));
  assign y1 = (-4'sd7);
  assign y2 = ((p11>=p1)*(5'd2 * p13));
  assign y3 = $signed(({3{(p6>=p17)}}<{(-$signed({1{(p14)}}))}));
  assign y4 = (&((~(-$signed({3{{2{(p6^p6)}}}})))));
  assign y5 = ((((b2>>>b4)&(|a1))!==$signed((~&{4{b3}})))>>>(+$unsigned({3{{4{p14}}}})));
  assign y6 = ((5'd2 * b0)?(a5===a4):(p11-b0));
  assign y7 = (a0==a4);
  assign y8 = (((p12<<p14)?$unsigned((p3==a3)):(b1===a5))||{4{(p10>>p4)}});
  assign y9 = ((~&a5)^~(b0-b4));
  assign y10 = (^(|$signed(p7)));
  assign y11 = (&(+a4));
  assign y12 = {1{(+{4{{1{(~{3{b3}})}}}})}};
  assign y13 = (~(p12>=p13));
  assign y14 = {2{p15}};
  assign y15 = (a2?b1:a1);
  assign y16 = (4'sd5);
  assign y17 = (~&((p6|p17)?(p0!=p1):(p5<=p13)));
endmodule
