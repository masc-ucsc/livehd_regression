module expression_00495(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd5)==((2'd1)<<(4'd9)))-((2'd1)?(-5'sd10):(5'd22)));
  localparam [4:0] p1 = ((-2'sd0)?(5'sd14):(2'd3));
  localparam [5:0] p2 = (2'sd0);
  localparam signed [3:0] p3 = {1{({2{((3'd0)||(4'd3))}}||{(2'sd0),{(5'd0),(2'sd0),(4'd6)},{2{(-5'sd11)}}})}};
  localparam signed [4:0] p4 = (^{(^(~(3'd6))),(^(~^(3'd5))),(&(+(-5'sd8)))});
  localparam signed [5:0] p5 = {{(4'd2),(3'd0),(3'sd1)},(~|(2'sd1))};
  localparam [3:0] p6 = (&({(((-4'sd4)^(2'd3))!={(4'd13),(3'd1),(3'sd1)})}&(&(~^{((-3'sd3)|(-3'sd0)),((5'sd8)>>(-3'sd3))}))));
  localparam [4:0] p7 = (2'd1);
  localparam [5:0] p8 = ({2{{(3'sd0),(5'sd0),(4'sd2)}}}?((-3'sd3)?(4'sd7):(5'd29)):(((2'd1)-(2'd3))|(3'd6)));
  localparam signed [3:0] p9 = {(5'd18),(5'sd4),(3'sd1)};
  localparam signed [4:0] p10 = ({4{(4'd11)}}>={3{(5'd21)}});
  localparam signed [5:0] p11 = {{(((2'sd1)<(5'd30))-((3'd4)<=(2'd0)))},{4{{4{(2'd2)}}}}};
  localparam [3:0] p12 = {(2'd0),(-4'sd5)};
  localparam [4:0] p13 = (2'd1);
  localparam [5:0] p14 = (-((~(4'sd5))>=(-3'sd3)));
  localparam signed [3:0] p15 = (((5'sd0)<<<(-4'sd4))<((-5'sd9)^~(-2'sd1)));
  localparam signed [4:0] p16 = ((+{1{{3{((-2'sd1)^~(3'd5))}}}})&&(~{(((4'd12)?(-5'sd5):(2'd1))?(+(2'd1)):((-5'sd11)?(5'd28):(2'sd0)))}));
  localparam signed [5:0] p17 = (|((~^(3'sd3))?(!(5'd28)):((-5'sd0)?(-3'sd1):(5'sd9))));

  assign y0 = ((3'd0)&((-5'sd15)!==(($unsigned({4{a0}})))));
  assign y1 = (|a5);
  assign y2 = {2{{2{(&a2)}}}};
  assign y3 = (+(+(^(a3==p1))));
  assign y4 = (b5!==a2);
  assign y5 = {3{b1}};
  assign y6 = (~(((p3^~p16)^~(&p14))>>>(4'd2 * {p2,p8})));
  assign y7 = (($signed(($signed(p6)+(p5)))&((p10||p4)>>>(5'd19)))==(3'sd3));
  assign y8 = {(p0?a3:a3),(a1?a4:p8),(-5'sd6)};
  assign y9 = (b5/p17);
  assign y10 = ((~|{{(p5<<p0),{p13},$signed(a4)}})>=((5'd28)===(&$unsigned((b2-a5)))));
  assign y11 = (^((+(~((~|a1)<<(~^b1))))^~(5'd2 * (^(a1!=a2)))));
  assign y12 = {3{(b5>>a4)}};
  assign y13 = (($signed($signed(($unsigned(a3)&$signed(b0)))))===((b1)?(a2):(b5*a3)));
  assign y14 = (&(4'sd6));
  assign y15 = (((a5?a4:a2)&&((p10^~a4)))+(((p6*a2)==(b5?p4:b4))&&$unsigned($signed((p5?a4:p2)))));
  assign y16 = $signed({2{{p8,a0,b5}}});
  assign y17 = {{((+{((b4?b0:a4)+{a1,a1,b3})})!=={(+(+(b3?a2:a0))),(!(a4?a5:b0))})}};
endmodule
