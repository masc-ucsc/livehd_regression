module expression_00439(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-((-5'sd6)===(4'sd5)));
  localparam [4:0] p1 = (|((3'sd2)<(-5'sd0)));
  localparam [5:0] p2 = ((-2'sd1)==(2'd1));
  localparam signed [3:0] p3 = ((3'd0)>>>{4{(4'sd0)}});
  localparam signed [4:0] p4 = {2{(~{(+(2'd0))})}};
  localparam signed [5:0] p5 = {3{(-3'sd3)}};
  localparam [3:0] p6 = {{(5'd0)},{({4{(3'd0)}}==={1{(5'sd9)}})}};
  localparam [4:0] p7 = ((!(5'd2 * (5'd25)))>>{(4'd13),(2'sd1)});
  localparam [5:0] p8 = {3{(-5'sd7)}};
  localparam signed [3:0] p9 = (((2'sd1)?(-5'sd1):(-5'sd2))===(4'd2 * (3'd2)));
  localparam signed [4:0] p10 = ((4'd14)?(3'd6):(-3'sd3));
  localparam signed [5:0] p11 = (3'd3);
  localparam [3:0] p12 = ({{({3{(-3'sd3)}}&(!(-(2'sd0))))}}!=(5'd2 * {(4'd6),(4'd7),(3'd4)}));
  localparam [4:0] p13 = (((~^((2'sd1)!=(3'd7)))<=((4'sd4)-(-3'sd0)))-(((5'sd8)%(2'd2))+((3'd5)%(2'd3))));
  localparam [5:0] p14 = (-((-2'sd0)<(-3'sd2)));
  localparam signed [3:0] p15 = (~(~&((^(5'd26))?(~(4'd14)):((3'sd0)?(4'd6):(4'sd4)))));
  localparam signed [4:0] p16 = (~&{(((-4'sd4)>(2'd1))^{4{(5'd10)}}),(-4'sd1)});
  localparam signed [5:0] p17 = (|(3'd7));

  assign y0 = (4'd14);
  assign y1 = (-((~(2'sd1))?(p5?a3:p15):(3'd2)));
  assign y2 = (+(p14?p11:b4));
  assign y3 = ({4{(a5>a0)}}>$signed(((a2?b5:b4)?{3{a2}}:{3{b4}})));
  assign y4 = (((p10>=a5)));
  assign y5 = (4'd2 * p8);
  assign y6 = ((~^(^{{p0,b4}}))?(3'd1):(^((2'sd0)^(~&b2))));
  assign y7 = (2'd1);
  assign y8 = {{{{(a3===b5)},{(b4<=b0)},((a3&&b2)==={b0,a5,a1})}}};
  assign y9 = {4{(!{2{p4}})}};
  assign y10 = {$signed($unsigned((!b1))),((a3==b5)^~{2{a1}}),{{2{b2}}}};
  assign y11 = {4{((b2?a2:p6)?(p8?p7:p4):(p6?b1:a5))}};
  assign y12 = ((&((!a2)>(p5<p7)))-{(p5==p7),$unsigned((p3^p6))});
  assign y13 = (~|{3{(p15?p1:b1)}});
  assign y14 = $unsigned((&(!({(b2^b4),(b0<<<a0),(a3^~b5)}))));
  assign y15 = (4'sd0);
  assign y16 = ({3{(!(+a5))}}<((&{2{b4}})<<<(b1?b3:a5)));
  assign y17 = (((p14&p1)?(b4?p3:p14):(p10-p15))<<<(((a1?b5:b0)^(a2===b3))<<((a1==p14)?(b2!=a0):(4'd2 * b2))));
endmodule
