module expression_00771(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^{3{{4{(3'd6)}}}});
  localparam [4:0] p1 = {1{(-3'sd1)}};
  localparam [5:0] p2 = {1{(-3'sd3)}};
  localparam signed [3:0] p3 = (!(~&{4{((2'd2)?(4'sd4):(-2'sd0))}}));
  localparam signed [4:0] p4 = (2'd3);
  localparam signed [5:0] p5 = (({(4'sd4),(-5'sd2)}>>>((2'd3)^(2'd1)))+(-({(2'sd1),(2'd2),(-2'sd1)}?{(3'd5)}:((-2'sd0)&(3'd0)))));
  localparam [3:0] p6 = (((5'sd15)?{(5'd17),(3'd1)}:{(5'd18)})>>(((2'sd0)?(-5'sd4):(5'd22))=={(4'sd2),(2'sd1)}));
  localparam [4:0] p7 = {4{(4'd12)}};
  localparam [5:0] p8 = (3'd0);
  localparam signed [3:0] p9 = (((-5'sd0)?(-4'sd5):(4'sd1))>>(~^(-5'sd3)));
  localparam signed [4:0] p10 = (4'sd2);
  localparam signed [5:0] p11 = ({{2{(4'sd3)}},{(3'sd1)}}>>>(((-4'sd4)+(-2'sd1))^~(~&(2'd2))));
  localparam [3:0] p12 = (((4'd12)>>>(2'd2))?{(2'd2),(4'sd6),(5'sd14)}:{(-5'sd11),(4'd2)});
  localparam [4:0] p13 = ((^{4{(2'd1)}})&((2'd0)<=(2'd0)));
  localparam [5:0] p14 = (2'd0);
  localparam signed [3:0] p15 = {4{(&{(4'sd0),(4'd12)})}};
  localparam signed [4:0] p16 = ((-5'sd1)?(4'd7):(4'd2));
  localparam signed [5:0] p17 = (6'd2 * ((3'd7)<=(2'd0)));

  assign y0 = (-(p6<<<p7));
  assign y1 = ((-((a2^a4)>=(b5!==a5)))-((3'sd2)?(5'd2 * p1):(a0?p14:b0)));
  assign y2 = ({(a3?a2:a5),{1{{2{a2}}}},{4{a3}}}==={4{{1{(a1?b5:b2)}}}});
  assign y3 = ((-{b4,b2,p13})<<{b5,b4});
  assign y4 = ({2{{3{a2}}}}>>>(p5?p1:b2));
  assign y5 = (p8-p1);
  assign y6 = ($unsigned((b3?b1:a0))!==(a3|a0));
  assign y7 = (~^(~|{3{{4{b2}}}}));
  assign y8 = $signed(((~&{(3'd1)})?($unsigned(a3)|(p1&p6)):({p12,p4}<=(b1?p1:a5))));
  assign y9 = (|(({1{p4}}^(p17?b3:a1))==({a3,a3,a0}|{3{b2}})));
  assign y10 = ((+((-5'sd8)+(2'd1)))^~($signed(b1)?(+p10):(a2)));
  assign y11 = (p15-p7);
  assign y12 = (((2'd1)?({1{a0}}?(2'd1):(p10?p17:p0)):((a5&&p6)^~(a4?p3:a4))));
  assign y13 = (({4{p1}}));
  assign y14 = (~|$signed((5'd2 * (a2>=p7))));
  assign y15 = (3'd3);
  assign y16 = {(((a1&p16)<$unsigned(b4))+($signed(p8)+{a1}))};
  assign y17 = {3{{2{b5}}}};
endmodule
