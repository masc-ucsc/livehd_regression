module expression_00025(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((3'd2)===(5'sd7))?((-3'sd2)?(3'sd3):(-3'sd3)):((-5'sd8)===(4'd2)))?(-2'sd1):((5'd2 * (3'd3))?{(3'd1),(3'd3)}:{(2'd2),(4'sd5)}));
  localparam [4:0] p1 = (((3'd1)?(4'sd1):(2'sd1))?{2{(3'sd1)}}:{2{(-5'sd14)}});
  localparam [5:0] p2 = ((5'd25)<<<(5'd17));
  localparam signed [3:0] p3 = {3{(4'd8)}};
  localparam signed [4:0] p4 = (|{3{(5'd2)}});
  localparam signed [5:0] p5 = (4'sd5);
  localparam [3:0] p6 = (((((2'd3)&&(-2'sd1))===((2'd1)<<<(2'sd0)))!=(((5'd1)||(5'd2))<=((3'd6)-(3'd5))))^~(((2'd2)<=(5'sd7))/(2'd2)));
  localparam [4:0] p7 = (~|(~&(~(-(((~&((5'd13)+(3'd4)))&((5'sd9)%(5'd20)))+(!(+(((3'd2)<<<(-4'sd0))+((4'd13)&(-5'sd5))))))))));
  localparam [5:0] p8 = ((+(5'd7))===(-4'sd3));
  localparam signed [3:0] p9 = (5'sd4);
  localparam signed [4:0] p10 = {(~|(3'sd1))};
  localparam signed [5:0] p11 = (&(((4'd14)?(3'd7):(2'sd1))^((3'd7)>(-4'sd7))));
  localparam [3:0] p12 = {2{(((2'd2)||(2'd3))<((3'd6)^~(2'd0)))}};
  localparam [4:0] p13 = (^{1{(+(~&(!(((4'd10)?(2'd2):(4'd10))?{2{(3'sd0)}}:(&(4'd9))))))}});
  localparam [5:0] p14 = {{{1{(3'd7)}},{2{(4'd7)}}},((5'd18)>={(4'd8),(5'd28),(4'd4)}),{((4'sd1)>(5'sd5)),{2{(-3'sd1)}},{2{(5'sd14)}}}};
  localparam signed [3:0] p15 = (-(&(~{{(2'd0),(2'sd1),(5'd12)}})));
  localparam signed [4:0] p16 = (~(3'sd1));
  localparam signed [5:0] p17 = ((3'sd1)?(((2'd1)<=(3'sd1))!==((5'd15)===(5'sd1))):(~((-2'sd0)&&(2'd3))));

  assign y0 = {4{b4}};
  assign y1 = ((3'sd0)-((3'd0)!=(2'd0)));
  assign y2 = (((b0===b1)+(~a3))!=((a0!=a3)^(a5<<p17)));
  assign y3 = {(4'd4),(|{{(^b5),{b5,a5}}})};
  assign y4 = (b1?a2:b1);
  assign y5 = (~{(((&a5)<={3{p16}})-(+(p16==p5))),(-(~&{3{{4{a4}}}}))});
  assign y6 = ((b5-p4)?(3'sd3):(p0>>b3));
  assign y7 = {(-2'sd0)};
  assign y8 = ({4{b5}}>(~|b5));
  assign y9 = {1{((^(p6?p7:b4))||$unsigned((~((p16>=p14)))))}};
  assign y10 = (~(p4||p13));
  assign y11 = ((~|p10)^~(|b1));
  assign y12 = (((a2|p9)<(p10&p13))+{(&({p15,p12}^~(p0>>>p9)))});
  assign y13 = ((((~|b2)>=(b1<<b1))===(|{$signed(b3)}))&{{3{p6}},(p1<<p17),(p12>=p1)});
  assign y14 = ((^(p16?p12:b0))?(b2&&p7):(p10?b4:b2));
  assign y15 = (5'd2);
  assign y16 = {(+$unsigned({(p2),(~p8)})),(-(~&(+(!({a5}))))),{$unsigned((~{($signed(p3))}))}};
  assign y17 = {4{p12}};
endmodule
