module expression_00931(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd1)>>>(-2'sd1))?((4'd2)?(2'sd0):(2'd1)):{1{(5'd30)}});
  localparam [4:0] p1 = {2{(((4'd11)>>>(5'sd5))>((-5'sd3)<<(3'd4)))}};
  localparam [5:0] p2 = ((-(((4'd6)^(5'd3))||(^(-(-4'sd6)))))>(|(((-3'sd3)?(4'd10):(3'd1))!=((4'sd4)&(3'd4)))));
  localparam signed [3:0] p3 = {1{{1{(&(((2'sd0)^(5'sd15))||{4{(5'd31)}}))}}}};
  localparam signed [4:0] p4 = {((-3'sd2)?(4'd9):(2'd3)),((2'sd1)?(-3'sd0):(5'sd13)),(|(-5'sd13))};
  localparam signed [5:0] p5 = (~(3'd0));
  localparam [3:0] p6 = (!((!(((5'd16)&&(5'd27))<=((-3'sd3)?(5'sd7):(5'd25))))+({(2'sd1),(2'd0),(4'sd4)}^~{(-3'sd3),(2'd3),(5'd7)})));
  localparam [4:0] p7 = (5'd2 * {2{(4'd14)}});
  localparam [5:0] p8 = ((^{4{(4'sd4)}})>(((2'd0)!==(3'd5))<<<((-4'sd3)^~(2'd1))));
  localparam signed [3:0] p9 = ((^(-((-2'sd0)?(-2'sd0):(-4'sd1))))?(^((~^(2'd3))^{4{(3'sd1)}})):((+(2'sd1))&&((2'd0)?(5'd9):(2'd2))));
  localparam signed [4:0] p10 = ((4'd13)>(-3'sd0));
  localparam signed [5:0] p11 = ((-5'sd15)>>(((3'd0)<<(5'sd9))&&{2{(5'd5)}}));
  localparam [3:0] p12 = ((~|((^(5'd5))<<<((3'd5)||(5'sd12))))?((+(2'sd0))?(^(3'sd3)):((-5'sd6)!==(-2'sd0))):(((3'd6)^(-2'sd1))>>{1{(5'd24)}}));
  localparam [4:0] p13 = {3{{3{(3'd7)}}}};
  localparam [5:0] p14 = ((4'd3)?(4'd1):(2'd3));
  localparam signed [3:0] p15 = ({4{(2'sd0)}}?{3{(2'd3)}}:((4'sd7)?(-3'sd2):(3'sd2)));
  localparam signed [4:0] p16 = ({(6'd2 * (5'd17))}&&(|((4'd15)|(4'd5))));
  localparam signed [5:0] p17 = ((&(4'd7))>>>({3{(2'd2)}}!=((4'sd0)<<(5'd18))));

  assign y0 = (3'sd2);
  assign y1 = (2'd1);
  assign y2 = (((4'd2 * a2)<<($signed(p17)))|({1{$signed(a5)}}=={4{b2}}));
  assign y3 = (~|{4{p14}});
  assign y4 = (5'sd0);
  assign y5 = ((2'd1)>=($unsigned($unsigned($signed(p9)))));
  assign y6 = (!(|((2'd3)/a0)));
  assign y7 = {4{(5'd7)}};
  assign y8 = $signed((2'd1));
  assign y9 = (~($signed(p17)?(p16?p12:p15):(~&p7)));
  assign y10 = (((p12?p3:p6)<$signed(p16))>>(((p11<<p6)>=(p2>=p9))));
  assign y11 = $signed(({2{{1{(~b5)}}}}!==$unsigned({3{{2{a4}}}})));
  assign y12 = (~&((((5'd2 * (~^(~^a2)))))|$signed(((p4!=p17)^((~|b1))))));
  assign y13 = {3{p6}};
  assign y14 = (^{3{$unsigned($signed(p8))}});
  assign y15 = (5'sd13);
  assign y16 = {b3,b3};
  assign y17 = (4'sd1);
endmodule
