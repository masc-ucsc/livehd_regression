module expression_00939(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{((-5'sd7)?(4'd5):(-3'sd1)),((4'd12)||(4'sd2))},{{2{((5'sd0)?(3'sd0):(2'sd1))}}}};
  localparam [4:0] p1 = {(~({((3'd1)?(2'd0):(-3'sd2))}?(~^(4'sd1)):(3'd5)))};
  localparam [5:0] p2 = (!(-((((2'd2)&(3'd1))/(-5'sd8))^~(~((~|(2'sd1))<(&(4'd9)))))));
  localparam signed [3:0] p3 = (~^(4'd2 * (4'd6)));
  localparam signed [4:0] p4 = ((~|{{(5'sd6),(3'd5),(5'd2)}})?((+(3'sd3))?(|(5'd18)):((4'd8)?(4'd7):(2'd1))):(~^(^{(4'd3),(3'sd1)})));
  localparam signed [5:0] p5 = (~^(&(-(&(&{2{(+(-2'sd0))}})))));
  localparam [3:0] p6 = {(-4'sd6)};
  localparam [4:0] p7 = ({(3'd2),(4'd12),(-5'sd0)}==(!(4'd10)));
  localparam [5:0] p8 = {1{{2{{3{{3{(-3'sd3)}}}}}}}};
  localparam signed [3:0] p9 = (&((((2'sd1)^~(5'sd14))+(6'd2 * (5'd17)))|((-{1{(5'd1)}})!=(&{(5'd3)}))));
  localparam signed [4:0] p10 = {((((5'd31)<(2'd0))!=={(5'd18),(-4'sd6),(5'sd10)})>=(^((~{(3'd4),(2'd3),(5'sd13)})||{(-3'sd2),(-3'sd1)})))};
  localparam signed [5:0] p11 = (((2'sd0)?(2'd2):(2'd0))?((-5'sd13)?(4'd2):(5'sd6)):((5'd28)?(3'd7):(3'd5)));
  localparam [3:0] p12 = {1{(5'd3)}};
  localparam [4:0] p13 = (2'd0);
  localparam [5:0] p14 = (-3'sd1);
  localparam signed [3:0] p15 = (2'd1);
  localparam signed [4:0] p16 = ((3'd5)?(-3'sd1):(5'd11));
  localparam signed [5:0] p17 = {3{(|(3'd5))}};

  assign y0 = ((((a2<=p12)>=(-a4))>=((b4||a1)>=(p13>>b0)))<<(((p17<<<p14)!=(b2===b1))>>((b4&b0)!==(a0!==a3))));
  assign y1 = (3'sd2);
  assign y2 = ({p14,b1,p16}==((b4>>b4)&(^b2)));
  assign y3 = $signed($unsigned({(p4==p16),(p15||a2)}));
  assign y4 = {({1{(4'd2 * p14)}}|{b2,p11,p15}),{{p12},{a0,p12,p8},(p14|p9)},(6'd2 * {4{p13}})};
  assign y5 = ((b5<=b3)?(a2<<<p12):(p17?a2:b3));
  assign y6 = (^((((!b1)=={3{a4}})==((b5>b1)!==(-b0)))==={4{(a4>=a1)}}));
  assign y7 = (~{2{(^(!(-((!b0)+(p5>a0)))))}});
  assign y8 = (2'd3);
  assign y9 = ((2'd1));
  assign y10 = ((2'd3)<(p4?a3:p0));
  assign y11 = ((a3===a1)<<<(p8?a2:p13));
  assign y12 = {3{((a1!==a3)&(+(!b0)))}};
  assign y13 = ($signed(($unsigned((!p4))?$unsigned((a2==p17)):$signed((p5>>a5)))));
  assign y14 = {4{(b1!=a0)}};
  assign y15 = ($unsigned(({2{b2}}>=(a4+a5)))!=(~^(~|({a3,a4}))));
  assign y16 = (!(3'd5));
  assign y17 = (((&(~|p0))^(p17<<p13))?((p4?p16:b2)||(p14|p9)):(&((p11+p12)<(&p12))));
endmodule
