module expression_00994(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&({((4'd9)|(-5'sd1)),((3'd4)<<<(4'sd0)),((5'd24)&&(2'd3))}+((~|{(4'sd0)})==(|(^(4'sd0))))));
  localparam [4:0] p1 = (5'd2 * (3'd0));
  localparam [5:0] p2 = (3'sd1);
  localparam signed [3:0] p3 = (~|((!(-{(!((-2'sd1)>>(4'd8)))}))|(((4'd5)&&(-3'sd3))+((4'd4)||(5'sd7)))));
  localparam signed [4:0] p4 = {(({(~^(-3'sd3))}<=((5'sd4)||(-2'sd0)))^(-{{{(4'd0),(2'd3),(3'd4)}},((4'sd6)^(-4'sd2))}))};
  localparam signed [5:0] p5 = ((2'sd1)-(5'sd3));
  localparam [3:0] p6 = (-{4{(+(4'd10))}});
  localparam [4:0] p7 = ((((-4'sd6)?(4'd11):(-3'sd0))<<((-2'sd1)?(3'd2):(4'sd4)))?(((5'd6)!=(4'd3))^((3'sd1)+(2'sd0))):((-(5'sd15))?(~(3'sd3)):((4'sd0)?(2'd1):(2'sd1))));
  localparam [5:0] p8 = ((3'd0)?(-2'sd1):(3'd3));
  localparam signed [3:0] p9 = {(({(-2'sd1),(5'sd12)}!=={(5'd1),(4'sd7)})<=(((3'd7)-(-4'sd4))>((3'd5)-(5'd18)))),{((5'd18)-(2'd2)),((-4'sd1)^(4'sd0)),{(5'sd15),(5'sd14)}}};
  localparam signed [4:0] p10 = ((((3'sd0)>>>(4'd11))||(~&(4'd10)))>=(-2'sd1));
  localparam signed [5:0] p11 = ({1{(2'sd1)}}?(~&(-5'sd2)):((4'd1)?(3'd4):(5'd3)));
  localparam [3:0] p12 = ((-5'sd11)|(5'd8));
  localparam [4:0] p13 = ((-4'sd7)^~(((2'd0)-(3'd5))===(5'sd9)));
  localparam [5:0] p14 = {(!{(2'd0)}),((-3'sd3)?(4'd2):(2'd1)),(-(~^(4'd12)))};
  localparam signed [3:0] p15 = (-((4'd3)?(-2'sd1):(3'sd2)));
  localparam signed [4:0] p16 = {2{(-2'sd0)}};
  localparam signed [5:0] p17 = (|(~&(((2'sd1)||(-3'sd2))?(~&(3'd6)):(^(-4'sd6)))));

  assign y0 = {3{{4{(3'd1)}}}};
  assign y1 = (-3'sd3);
  assign y2 = (~|$unsigned({{b2,p15},(p13?b2:a2),$unsigned(b1)}));
  assign y3 = $unsigned((~|{4{(b1>=p15)}}));
  assign y4 = (2'd3);
  assign y5 = ((4'd4)?(3'd0):(b4==b4));
  assign y6 = {(a4?p6:a1),((p14<=a3)|{p10,b0}),((a0>b4))};
  assign y7 = (p17&&p17);
  assign y8 = $unsigned((($signed(a5)?(p0&a3):{3{b5}})?({3{p14}}?(b4<<b4):{3{b4}}):{2{(p15^a2)}}));
  assign y9 = ({((a2<<p12)?(a4?b0:p1):(~&b3))}>{(~p11),(b0?p0:b0),(~|a0)});
  assign y10 = ((-((b2!==a0)>>(b2+p0)))=={{(p8+p6),(~|p7)}});
  assign y11 = (b2<b4);
  assign y12 = (~|(((+(+a0))||(b4?p0:p6))>>((a0===a2)^~(p3>>>a4))));
  assign y13 = ({({b1}===(4'd14))}-{{p12,a2},(4'd2 * b0)});
  assign y14 = ((((p8^p0)==(a2^~p11))>{3{p1}})>>({1{(p10&p3)}}<((p11>>>p4)<{4{p5}})));
  assign y15 = (((b5===a4)+(p4-p4))==((a4!==a1)===(b2>=a5)));
  assign y16 = (3'sd3);
  assign y17 = ({4{p12}}&({4{p10}}>>>(~&p0)));
endmodule
