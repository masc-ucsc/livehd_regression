module expression_00008(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{3{(3'd3)}}}};
  localparam [4:0] p1 = (-{((2'd2)?(3'd6):(-5'sd2))});
  localparam [5:0] p2 = {{(3'd6)},((4'sd2)>=(5'd9))};
  localparam signed [3:0] p3 = ((((5'd21)>>>(4'd14))?((4'd10)/(3'd0)):((2'd2)%(4'd12)))&&(((4'd12)?(5'd26):(4'sd6))|((-2'sd1)==(5'd13))));
  localparam signed [4:0] p4 = (5'd0);
  localparam signed [5:0] p5 = (^{((((5'sd14)&(5'd0))>(~&{(4'sd2)}))!==(&((^((-3'sd2)&&(-4'sd5)))===(^((2'd1)||(2'sd0))))))});
  localparam [3:0] p6 = ((5'd23)?(2'sd0):(2'sd0));
  localparam [4:0] p7 = ({{(-2'sd1),(-3'sd1),(2'd1)},(~(3'd3)),((-3'sd0)^(3'd7))}>>>{((2'd1)^(5'd28)),((-5'sd5)?(5'd12):(5'sd6)),{4{(3'sd2)}}});
  localparam [5:0] p8 = ({(-5'sd14),(4'd13),(5'd17)}!={(3'sd0),(4'sd2),(-3'sd1)});
  localparam signed [3:0] p9 = {4{({4{(5'd14)}}<=((2'sd1)>(2'sd0)))}};
  localparam signed [4:0] p10 = (5'd2 * ((2'd3)&(5'd8)));
  localparam signed [5:0] p11 = ((((4'd6)^~(4'd11))<<(+(3'd1)))<(~&((4'd12)&(5'd21))));
  localparam [3:0] p12 = (~&(&(^(~^(5'sd1)))));
  localparam [4:0] p13 = {4{{2{(3'd0)}}}};
  localparam [5:0] p14 = {((5'd19)?(4'd15):(5'd6)),((2'd1)?(5'd28):(4'd2)),(6'd2 * (5'd3))};
  localparam signed [3:0] p15 = {(2'sd0)};
  localparam signed [4:0] p16 = (((2'd3)?(4'sd0):(3'd4))==(3'd6));
  localparam signed [5:0] p17 = {({(3'd2),(3'sd1)}+(~|{(3'd4),(4'd0),(4'd12)}))};

  assign y0 = (^(~|$signed($signed({(&{4{a3}})}))));
  assign y1 = (|($unsigned((+p10))/b1));
  assign y2 = (|(((|((|b5)^(a0<<a0)))===$unsigned(({a5}!=(-b1))))>{(((~&b3)!==(!a2))<<<({p1,p15,p1}>(~p9)))}));
  assign y3 = (4'd3);
  assign y4 = {(({b5,a1}&&(a1>=a4))===((b3==b4)+(b2==b5)))};
  assign y5 = (2'sd0);
  assign y6 = (-5'sd6);
  assign y7 = (-((&(a0?a1:b2))?$signed(((~&(b3?a2:b3)))):(~|(-(b4?b4:a3)))));
  assign y8 = ({1{((b2^~a4)^(b1-p0))}}?{4{a1}}:((b4!==a2)||(b3<<<a2)));
  assign y9 = {2{{2{(!(|(4'sd5)))}}}};
  assign y10 = {{{1{(b5?b1:b2)}},{3{a0}}},{1{({b0,b5}?(b3?b3:a0):{a5})}},{({2{p10}}?(a1?b4:a4):(a0?a0:a1))}};
  assign y11 = {{p14,p10,p15},$signed((-3'sd3))};
  assign y12 = (((~&a1)>>>(p1^p13))>=(|(4'd2 * (b1===a0))));
  assign y13 = (((3'sd0)>=(-(~^(~^(a0+a4)))))===(+{(5'sd12),(-5'sd5),(a0||a0)}));
  assign y14 = (&{(-(!(5'd12)))});
  assign y15 = {(((p15<<<a2)|{a1,p17})<((~|(b1&b4))!==(-2'sd1)))};
  assign y16 = $unsigned(((p17?b5:a1)?{3{p5}}:{3{p7}}));
  assign y17 = (4'sd3);
endmodule
