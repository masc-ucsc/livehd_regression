module expression_00196(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd4);
  localparam [4:0] p1 = (5'd2 * {(2'd0),(2'd0)});
  localparam [5:0] p2 = ((&(2'd2))?(~(5'sd7)):((3'd3)+(5'sd3)));
  localparam signed [3:0] p3 = ({((3'd2)>=(2'd0)),((5'd5)?(4'sd6):(-5'sd12))}>>(5'sd8));
  localparam signed [4:0] p4 = (~((4'd0)<<(2'd1)));
  localparam signed [5:0] p5 = {(^{3{(4'd2)}})};
  localparam [3:0] p6 = {{(2'd0),(4'd14),(4'd4)},((~&(2'd1))&&((4'd7)-(2'd1))),(((-5'sd11)^(5'd17))>>{(5'sd9),(2'd3),(3'sd2)})};
  localparam [4:0] p7 = (~{4{{2{(5'd30)}}}});
  localparam [5:0] p8 = (|(2'd1));
  localparam signed [3:0] p9 = (|(({(3'd3),(3'd0),(5'd24)}&{(5'sd1)})^~(((5'd6)+(4'd13))===(^(5'd18)))));
  localparam signed [4:0] p10 = {{(|(((3'd1)|(2'd2))?{(-4'sd6),(-4'sd2),(-2'sd1)}:((2'd3)?(4'sd3):(-5'sd4)))),(((4'd2)===(-3'sd1))?{(4'd5),(5'd21)}:(+(-4'sd4)))}};
  localparam signed [5:0] p11 = ((3'd3)%(3'd6));
  localparam [3:0] p12 = {2{(2'sd1)}};
  localparam [4:0] p13 = (|{4{(2'sd0)}});
  localparam [5:0] p14 = (2'sd0);
  localparam signed [3:0] p15 = (|((((-4'sd2)?(5'sd3):(-5'sd14))>>>((5'd4)?(-2'sd1):(4'd12)))+(~|(((3'd0)<<<(2'd3))===((4'd2)?(4'd13):(-5'sd7))))));
  localparam signed [4:0] p16 = ((&((2'd3)?(5'd26):(-5'sd9)))?((-5'sd0)?(4'sd7):(3'd3)):((5'd9)?(5'd29):(5'd18)));
  localparam signed [5:0] p17 = ((2'd3)+((2'sd0)>>(2'sd0)));

  assign y0 = ({((p16|p10)<{p12,p4,p7}),((a0!=p2)<<{p10,p4,p7})}<={(p8<<<p0),(p10>=p2),(p17^p8)});
  assign y1 = ({4{a0}}?(4'sd3):({3{b4}}?(p14>b1):(b2?b5:a4)));
  assign y2 = (((p9>=p4)>>(p0||p11))&{2{(p6>>p3)}});
  assign y3 = {2{(~|({a2,p10,p3}^~(!p2)))}};
  assign y4 = (|(((b3<p10)|{3{p5}})>>>(^(+(-{3{p10}})))));
  assign y5 = ((!p7)?{2{p9}}:(p12>>p4));
  assign y6 = {a2,b2};
  assign y7 = {(6'd2 * p7),(2'd2),(3'd4)};
  assign y8 = (b2?a4:a5);
  assign y9 = (2'sd0);
  assign y10 = (~^((~^(-4'sd3))==={(-2'sd1),$unsigned(b2)}));
  assign y11 = {3{{p0,p14,a4}}};
  assign y12 = (|p5);
  assign y13 = (~(~(^((p13^b0)<(~(p16>>a4))))));
  assign y14 = ($signed((4'sd5))&{4{b1}});
  assign y15 = {3{$signed({3{(3'sd2)}})}};
  assign y16 = {((b3^a4)!==(b5>a0)),({2{a3}}>>{4{p13}})};
  assign y17 = ($signed((2'sd0)));
endmodule
