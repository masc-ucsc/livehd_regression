module expression_00977(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({{(4'd11),(4'd10),(4'd11)}}?(^(&(2'sd0))):{(^(5'sd12))});
  localparam [4:0] p1 = ((!((^{4{(5'sd3)}})<<((-2'sd0)-(2'sd1))))+{2{{((5'sd3)-(2'd2))}}});
  localparam [5:0] p2 = ((|{3{(2'd2)}})<<((5'd26)>>>(3'sd1)));
  localparam signed [3:0] p3 = {({(2'd2),(5'd30)}?(|(5'd12)):(+(2'd2))),{(4'sd5),(|(4'sd6)),{(2'd2),(2'd3),(-3'sd1)}}};
  localparam signed [4:0] p4 = (~|(&(3'd0)));
  localparam signed [5:0] p5 = (!(3'd0));
  localparam [3:0] p6 = (~(+(~^(~^((3'd2)&(3'd0))))));
  localparam [4:0] p7 = ((3'd3)>(2'd0));
  localparam [5:0] p8 = (~|{2{{{4{(4'sd4)}}}}});
  localparam signed [3:0] p9 = (~&(3'sd3));
  localparam signed [4:0] p10 = (~|(4'd6));
  localparam signed [5:0] p11 = ((2'sd1)?(4'sd4):(2'sd1));
  localparam [3:0] p12 = (2'sd1);
  localparam [4:0] p13 = ((-5'sd8)>=(3'd6));
  localparam [5:0] p14 = ({3{(-4'sd0)}}?(&{4{(5'd17)}}):((3'd3)^~(-4'sd4)));
  localparam signed [3:0] p15 = (~^{(&(~|({(5'd18),(5'd30)}?((3'sd1)?(2'd1):(-3'sd1)):{(5'd4),(2'sd0)}))),(&(((3'd4)?(-3'sd3):(2'd1))^~(&((4'sd3)<<<(-5'sd2)))))});
  localparam signed [4:0] p16 = ({4{(4'sd3)}}^~{1{{(-4'sd5),(2'd2),(2'd0)}}});
  localparam signed [5:0] p17 = {3{(4'd4)}};

  assign y0 = ((b5?a3:b2)?(|b0):(!b3));
  assign y1 = ((p13<p12)<={2{p14}});
  assign y2 = (~^{(4'd2 * p0),(p2<=p3),(~|a5)});
  assign y3 = {(~&{{{p0,p11,p8},(^{p4,p14})}})};
  assign y4 = {4{(b5>>>a5)}};
  assign y5 = ($signed((5'd10))===((b1)));
  assign y6 = ((4'd11)<=$unsigned(({4{p11}}!=(p6^~p9))));
  assign y7 = (+(-(~&(p7>b0))));
  assign y8 = (~|((+(~&b4))/p9));
  assign y9 = ({(p3!=p9),(b0===b4),{p10,p2}}<=(((b4)&$unsigned(b4))<<((b5<<<a2)===$unsigned(a3))));
  assign y10 = {3{{1{{{a0,b2,a5},(~^p11),(^a0)}}}}};
  assign y11 = ((~|(~{2{p3}}))?(-(~(p7?a3:a3))):{1{(&(&{3{b2}}))}});
  assign y12 = ($unsigned(b0)<=(p3!=p13));
  assign y13 = (~^(4'd2 * (^(5'd27))));
  assign y14 = {p13,p13,a1};
  assign y15 = (({3{a5}}+(b5<<a0))^~{2{(b4<<p14)}});
  assign y16 = (({3{a3}}==={4{a4}})<<({1{{1{a4}}}}&(p15||p15)));
  assign y17 = ({4{{1{$unsigned({2{a0}})}}}});
endmodule
