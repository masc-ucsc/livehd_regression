module expression_00273(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(((5'sd9)||(-4'sd2))^(2'sd1)),{(((4'd0)!==(4'd3))^~{(3'd1),(2'd0)})}};
  localparam [4:0] p1 = (^((((4'sd1)>>>(5'd26))<<<{(2'd2),(-5'sd15)})==(-{(3'sd0),(-4'sd4),(3'd7)})));
  localparam [5:0] p2 = (((4'd2 * (4'd8))<<((5'd7)?(5'd0):(5'd14)))^(((4'd8)?(5'sd15):(3'd3))===((3'd1)>>(3'sd3))));
  localparam signed [3:0] p3 = (~^(-(~(+((2'd0)==(3'd0))))));
  localparam signed [4:0] p4 = (|(-5'sd2));
  localparam signed [5:0] p5 = ((2'sd1)?(3'd2):(2'sd0));
  localparam [3:0] p6 = (~^(4'sd6));
  localparam [4:0] p7 = (!(((-4'sd3)>=(-4'sd0))>=(+(~^(3'sd0)))));
  localparam [5:0] p8 = ((~^(((4'd6)?(-3'sd3):(3'd2))>(~^((4'd6)&(3'd5)))))&(+(|(~&(~&((-2'sd0)<(2'd3)))))));
  localparam signed [3:0] p9 = (-5'sd12);
  localparam signed [4:0] p10 = ((((-4'sd0)?(5'd14):(3'd0))>>{(-2'sd0)})?(-3'sd0):(((-3'sd3)?(3'd5):(-4'sd4))===(-4'sd0)));
  localparam signed [5:0] p11 = ((^(~(3'd6)))?{4{(-4'sd5)}}:{2{(5'd7)}});
  localparam [3:0] p12 = (~|(~((~&(4'd5))<<((-3'sd0)^~(2'd3)))));
  localparam [4:0] p13 = {((~&(2'sd1))<<<(~|(4'd0))),{1{((3'd2)===(2'd2))}}};
  localparam [5:0] p14 = ((5'd26)|(-4'sd4));
  localparam signed [3:0] p15 = (-((~(4'd4))?((5'sd8)!==(5'd25)):((4'sd7)^(-2'sd1))));
  localparam signed [4:0] p16 = (^(|(((^(3'd2))|(-5'sd9))|((-(3'd3))?((2'd0)?(2'sd1):(5'd31)):((3'd5)|(5'd12))))));
  localparam signed [5:0] p17 = (2'd0);

  assign y0 = ({4{{3{p5}}}}<=({1{(b1===b2)}}<<{1{(p13>>>p5)}}));
  assign y1 = $signed((4'd8));
  assign y2 = {{(p3?p11:p6)},((2'd0)?(a4===a2):(p16<<p4)),((p0?p1:p9)?(-5'sd11):(6'd2 * p13))};
  assign y3 = ((a2?a2:p3)?(a1!==b5):(3'd5));
  assign y4 = {2{(p13|b1)}};
  assign y5 = (|{2{(+((a2&p3)?{p9,p10}:{3{b2}}))}});
  assign y6 = $unsigned(p6);
  assign y7 = {2{(-(~|(^{2{b3}})))}};
  assign y8 = ((((a3||a3)||(a3<<b5))==={(b3<=b1),(~|b3),(b2?a0:a0)})<<(({4{p6}}?(4'd2 * b0):{p16,p5,a3})+((a5^p13)>(p4>=b5))));
  assign y9 = (6'd2 * (3'd1));
  assign y10 = (3'sd3);
  assign y11 = (^((((~|b2))>>(b5&b3))==((b5>>>b3)!==(a4>=b0))));
  assign y12 = (2'd3);
  assign y13 = (~&(a2?b5:a4));
  assign y14 = (({2{p4}}?{1{p5}}:{p2})!=(-3'sd0));
  assign y15 = ((-2'sd0)===$signed({a2}));
  assign y16 = ((6'd2 * b2)/a3);
  assign y17 = {4{{2{b5}}}};
endmodule
