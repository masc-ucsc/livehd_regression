module expression_00777(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((&(3'sd2))?((-2'sd0)===(2'd3)):((5'd11)&&(5'd20)));
  localparam [4:0] p1 = (((2'd1)||(-5'sd8))<((-5'sd6)?(-5'sd12):(-3'sd3)));
  localparam [5:0] p2 = {4{(~&((3'd5)?(2'd1):(4'd12)))}};
  localparam signed [3:0] p3 = ((|(-4'sd2))+((|((5'sd15)?(3'd5):(2'sd0)))!==(5'sd11)));
  localparam signed [4:0] p4 = (((-2'sd0)-(2'd0))!=={1{(3'd2)}});
  localparam signed [5:0] p5 = (((3'd2)?(4'sd1):(3'd0))?(-4'sd6):((2'd1)?(-3'sd3):(-4'sd5)));
  localparam [3:0] p6 = ((~(-2'sd0))>=(~|(3'sd2)));
  localparam [4:0] p7 = ((&{1{{2{(4'd11)}}}})?(-(~^(~|(-4'sd2)))):(|((3'sd2)?(2'sd0):(5'd22))));
  localparam [5:0] p8 = (+(+(-4'sd7)));
  localparam signed [3:0] p9 = {((3'd5)&&(4'sd4)),{(5'sd3),(-5'sd0),(5'd14)}};
  localparam signed [4:0] p10 = {2{(-(5'd2 * {4{(5'd18)}}))}};
  localparam signed [5:0] p11 = {(-4'sd3),((5'd6)<(4'd9)),{(2'sd0),(4'd2),(3'd2)}};
  localparam [3:0] p12 = (4'd2 * ((2'd3)|(2'd3)));
  localparam [4:0] p13 = {{(5'd10),(2'sd0),(3'd3)},((-5'sd15)!==((-3'sd1)>>>(-5'sd5))),(-2'sd0)};
  localparam [5:0] p14 = ((((4'd2)<<(-5'sd14))==((2'd2)<=(4'd15)))<={3{(6'd2 * (4'd13))}});
  localparam signed [3:0] p15 = ((+{{(5'd24)}})?(^((-5'sd3)&&(-3'sd3))):(-5'sd0));
  localparam signed [4:0] p16 = {{(2'd1)},(3'sd2)};
  localparam signed [5:0] p17 = (((4'd3)?(4'd13):(2'd0))&(5'd2 * ((2'd2)>>>(4'd3))));

  assign y0 = (~^$unsigned(((|(^($signed(p17)?(~^p4):$unsigned(p8))))-($signed($unsigned(p14))>>(p9?p8:p16)))));
  assign y1 = (2'd1);
  assign y2 = $unsigned(({(p16+p17)}>=$signed((p6+p9))));
  assign y3 = ((((p16+p15)-(p4|b4))>((p11^~p15)^~(p5?p14:a0)))>=(((p16-p5)&&(p2?a0:p10))^~((p13<=p10)&&(p1<<p17))));
  assign y4 = $unsigned(((~|(((p17<=p11)==(b4!==b5))))==(~$unsigned(($unsigned(p3)<=(b4!==b4))))));
  assign y5 = ({(a5<b3),(&b5),(&b4)}?(!(+(b2?a2:a0))):((a5===b2)||{b3}));
  assign y6 = (4'd13);
  assign y7 = {(({p5,b1,a2}-(b2?a4:p11))!=(&(p8&&a1)))};
  assign y8 = (&(~^(~^{{(~^(|(&(~^{p8}))))},{{p1,p12},(^p12),(+a5)}})));
  assign y9 = (~|((~^(~^($unsigned((p3&&p0))||$signed((a0)))))||(((!b3)===(-a1))===(!(-$signed(b3))))));
  assign y10 = ((|(&((b5>b5)!==(-5'sd0))))&(2'd3));
  assign y11 = (!(+(3'd0)));
  assign y12 = ({{p12,a4,b3}}?{3{a4}}:{{3{p7}}});
  assign y13 = {((p14==p7)>=(p10>>p5)),(5'd2 * (^p6))};
  assign y14 = (~(^((~|{{3{b0}},{4{p0}},(-b2)})>>>(|((p6?b0:p0)^~{3{a3}})))));
  assign y15 = (-3'sd0);
  assign y16 = (a0<<a2);
  assign y17 = {(|p13),(a4!==a4)};
endmodule
