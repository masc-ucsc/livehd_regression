module expression_00152(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (4'sd7);
  localparam [4:0] p1 = (2'd0);
  localparam [5:0] p2 = {{(~(~(3'd3)))},(+(~(~&(3'sd2)))),({(2'd2)}<<{(2'sd0),(4'd12)})};
  localparam signed [3:0] p3 = (^(((3'd7)<<<(5'd24))>=((4'd1)^(2'd1))));
  localparam signed [4:0] p4 = (5'd2 * ((3'd6)||(3'd2)));
  localparam signed [5:0] p5 = (&{((-(2'd0))?{(2'd2),(3'sd3)}:((4'sd7)<(5'd28))),(~&{(-5'sd13)})});
  localparam [3:0] p6 = ({{4{(-5'sd13)}},(5'd15)}?{(2'sd0),{(4'd3),(5'sd12)},{(-2'sd1)}}:{{{(5'd6),(2'd0)}}});
  localparam [4:0] p7 = ({3{((2'd3)>>(5'sd4))}}-(((-5'sd9)^(4'd9))|((3'sd2)-(5'd17))));
  localparam [5:0] p8 = ((5'd11)===((-3'sd1)|{4{(2'd1)}}));
  localparam signed [3:0] p9 = ((~^(|((2'sd0)<(4'd15))))?({(3'sd1),(5'sd13),(4'sd6)}&((-3'sd3)<=(2'd2))):({2{(-3'sd1)}}>>{(5'sd10),(5'd10),(3'sd0)}));
  localparam signed [4:0] p10 = ((~^((+(~(-5'sd8)))<<<{4{(5'd15)}}))>>(((4'sd4)>=(4'sd2))>>>(+((2'd1)^~(3'sd2)))));
  localparam signed [5:0] p11 = (({1{(-2'sd0)}}?(-(4'd5)):{2{(5'd1)}})==((~&((3'sd3)?(5'd7):(4'sd1)))>>>(~^((2'sd1)==(2'd1)))));
  localparam [3:0] p12 = (-5'sd2);
  localparam [4:0] p13 = ((~&{(5'd12)})^{(((4'd14)===(4'd2))!=={3{(-2'sd0)}})});
  localparam [5:0] p14 = (4'sd0);
  localparam signed [3:0] p15 = (+{2{{((5'd17)-(4'sd0))}}});
  localparam signed [4:0] p16 = (3'sd1);
  localparam signed [5:0] p17 = {3{{2{(-2'sd1)}}}};

  assign y0 = $unsigned((+((a0*a0)===(a4!==a0))));
  assign y1 = {4{{4{a1}}}};
  assign y2 = ($signed($unsigned({4{{3{a5}}}}))&(2'd0));
  assign y3 = (p2>=p12);
  assign y4 = {{{{3{(a0?p2:b5)}},((p17!=b4)&(p10>>>p0))},{1{({2{(b3<=a3)}}!=={a0,b2,a3})}}}};
  assign y5 = (-{(((b1>>p6)^~{(~&p16)})>>(-{(^{p0,p1,p4}),(a1===b3)}))});
  assign y6 = (3'sd1);
  assign y7 = (p2?b5:p4);
  assign y8 = ((a2?a0:b3)?({1{(b5<p6)}}):{2{(b1>>b3)}});
  assign y9 = ((!p1)?(~^b0):(p4?a2:p3));
  assign y10 = ((p2?b1:b5)?(b1^b5):(!(~&p17)));
  assign y11 = ((-p15)>(p13!=p2));
  assign y12 = ((a2^~b0)?(4'd2 * a0):(b0+a2));
  assign y13 = (^(-(~|(((&p8)?(&a3):{p15})?({4{b2}}>>(b1<=p1)):((b3?a1:p8)<=(~&a4))))));
  assign y14 = (~|(((-(p3!=b2))/p7)^((4'd7)==(~p11))));
  assign y15 = ((((p2|p11)^~(4'd2 * p8))&((a4!==a4)>>{3{p4}}))==(((p15?p2:p4)>(p17<b3))>{p14,p16,p12}));
  assign y16 = ((&((p9+p7)<=(4'd8)))||(|{4{{p17,p9}}}));
  assign y17 = ({3{a3}}+((b3>p10)<={3{p13}}));
endmodule
