module expression_00200(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{{((2'sd0)?(-4'sd2):(-4'sd6))},((-2'sd0)-(4'sd0)),((3'd0)?(-4'sd7):(5'sd6))}};
  localparam [4:0] p1 = ((-5'sd14)^(3'd3));
  localparam [5:0] p2 = (|(^{1{(~(~&{4{(4'd2)}}))}}));
  localparam signed [3:0] p3 = ((&((4'sd7)&&(2'd2)))?((-(-4'sd1))!==((3'sd3)-(2'sd1))):(2'sd1));
  localparam signed [4:0] p4 = (((3'd7)^~(3'd6))==(5'd2 * (3'd5)));
  localparam signed [5:0] p5 = (((2'd2)-((4'd9)<<(-5'sd5)))<<(((5'd1)?(5'd2):(3'sd2))&(3'd5)));
  localparam [3:0] p6 = {2{(&{2{{3{(-2'sd0)}}}})}};
  localparam [4:0] p7 = ({2{(5'd9)}}^{(3'd0)});
  localparam [5:0] p8 = (&((3'sd0)-(3'd1)));
  localparam signed [3:0] p9 = ((2'd0)?((5'd2)%(4'd6)):(4'sd5));
  localparam signed [4:0] p10 = (((4'd14)<<(-2'sd0))^{(2'd2)});
  localparam signed [5:0] p11 = {{{{(5'd13)},{4{(4'd5)}},((5'sd2)+(3'd1))}}};
  localparam [3:0] p12 = (2'd0);
  localparam [4:0] p13 = (((4'd1)-(3'sd3))*(3'd6));
  localparam [5:0] p14 = ((|{(3'd2),(5'd31),(5'sd15)})>({(5'sd7)}<<(^(-5'sd10))));
  localparam signed [3:0] p15 = (~|((-4'sd6)?(3'd4):(4'sd6)));
  localparam signed [4:0] p16 = (-(-(~(2'd2))));
  localparam signed [5:0] p17 = ({({2{(-4'sd7)}}&&((2'd0)<(2'd0)))}&&{1{({(-5'sd0)}&&((5'd12)&(2'sd1)))}});

  assign y0 = {($unsigned($unsigned(($signed((~&((p6>p14)^~(b5<a3)))))))<<(3'sd3))};
  assign y1 = (&{p14,b3,p4});
  assign y2 = (~^(^(({a0}>{b3,b2})!=={b1,a2,b0})));
  assign y3 = {{a0},(b0?p12:a3)};
  assign y4 = (5'd12);
  assign y5 = $signed($signed((((p7>>p12)!=(5'd14))<<<((5'd28)!=$signed((~&p6))))));
  assign y6 = (+(+$signed($signed(({(2'd0)}<(^({2{b5}}<=(5'd31))))))));
  assign y7 = (!(+{3{{{3{(^p9)}}}}}));
  assign y8 = (((p14>>p1)<<<(p9>=p5))&({p9,p4,p16}|(a1&p14)));
  assign y9 = {4{(~^a2)}};
  assign y10 = (&(2'sd0));
  assign y11 = (((p13<<<a4)%b1)!=((p13/p15)*(p5>>a4)));
  assign y12 = (-2'sd1);
  assign y13 = ((+$signed(p8)));
  assign y14 = ((p2&p17)?(p15?p6:p10):(a0&&p13));
  assign y15 = ((4'd5)?(p4?p6:p11):(|(3'sd0)));
  assign y16 = {2{((5'd2 * a0)!==(^b4))}};
  assign y17 = ((3'sd3)+(^(a0|a4)));
endmodule
