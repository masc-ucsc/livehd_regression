module expression_00302(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{(3'sd1)}};
  localparam [4:0] p1 = (6'd2 * ((5'd6)===(4'd11)));
  localparam [5:0] p2 = {(^(4'sd4)),(-(-3'sd0)),((3'sd0)^~(3'd0))};
  localparam signed [3:0] p3 = ((4'd5)===(2'd3));
  localparam signed [4:0] p4 = (2'sd0);
  localparam signed [5:0] p5 = {{4{(4'd1)}},(((-5'sd1)||(-4'sd5))&(&(-2'sd1))),{(-2'sd1),(-2'sd1),(-5'sd3)}};
  localparam [3:0] p6 = (((&(-4'sd5))>>>((5'sd3)>>(4'sd6)))>{(4'sd4),(-2'sd1),(4'd15)});
  localparam [4:0] p7 = (~^(~|(~^(((2'sd1)?(3'd7):(3'sd0))?(!{{(4'd0),(2'sd1),(3'd7)}}):(4'd8)))));
  localparam [5:0] p8 = {1{{{((2'd2)>>(4'd15)),((4'd9)^(2'd3)),{4{(5'd19)}}}}}};
  localparam signed [3:0] p9 = ((((2'd3)===(2'd1))?((-5'sd7)^~(3'sd2)):(~^(3'd4)))&&(((5'd15)|(-3'sd2))?(4'd2 * (2'd3)):(~|(2'sd1))));
  localparam signed [4:0] p10 = (^(2'sd1));
  localparam signed [5:0] p11 = (~&(5'd14));
  localparam [3:0] p12 = (^((((-3'sd3)>>>(-4'sd2))>((2'd1)<<<(3'd0)))>({4{(4'd0)}}!==((2'sd1)^(-2'sd1)))));
  localparam [4:0] p13 = {2{(-2'sd1)}};
  localparam [5:0] p14 = ((4'sd7)?(3'sd0):(-4'sd0));
  localparam signed [3:0] p15 = ((((5'sd9)|(3'd0))^((-3'sd1)?(2'sd1):(3'd5)))<(((2'sd1)&&(3'sd3))>>((-2'sd1)||(3'd6))));
  localparam signed [4:0] p16 = {(&(~(((5'd0)-(5'd7))|(4'sd7))))};
  localparam signed [5:0] p17 = (~^(((~|(5'd27))==={(4'sd4),(-4'sd5),(5'd8)})>=((~&(2'sd1))&&{(5'sd14)})));

  assign y0 = $signed({2{{4{p15}}}});
  assign y1 = (b3<<<p8);
  assign y2 = ((+{4{p14}})?{1{((~&p9)?(p1|p2):(a1?p3:p5))}}:((~|p0)?$unsigned(p10):(-b2)));
  assign y3 = (-4'sd4);
  assign y4 = {4{((a2?a1:b3)===(b2?b4:b3))}};
  assign y5 = ({3{p3}}+(5'd8));
  assign y6 = ((b1?a2:a4)?(5'd2 * b1):(b1?b1:b2));
  assign y7 = {(^(a4==b2)),(a5>=b5),(p0&&a5)};
  assign y8 = (+({(2'd1),({3{{1{p17}}}}),{4{(^a1)}}}));
  assign y9 = {4{($signed(p7)<<<(a4>>p1))}};
  assign y10 = (^(((-2'sd1)<<{1{p8}})<<<(2'd0)));
  assign y11 = (({1{b3}}?(a5>>a1):{b4,a3,a0})|{{3{a0}}});
  assign y12 = (((b5>b5)+(5'd6))&(-4'sd1));
  assign y13 = ({1{((p16&&p1)|(~|{2{p0}}))}}<=((p8>>>p13)^~(p13>>>p7)));
  assign y14 = (((a1?p0:a0)&&({a1,b5,a1}<<(!p10)))==((~&(p5+a0))?{2{a2}}:$unsigned((b0<<<a0))));
  assign y15 = (+(~(-2'sd0)));
  assign y16 = ((^(b3+b1))%b0);
  assign y17 = {b0,p14};
endmodule
