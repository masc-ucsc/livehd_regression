module expression_00165(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~(4'd3));
  localparam [4:0] p1 = ({((-4'sd6)?(2'd3):(4'd9))}?((2'sd1)?(3'd3):(-4'sd6)):{(3'd3),(-2'sd1)});
  localparam [5:0] p2 = (-(&(+((-(+((-3'sd2)?(2'd0):(5'sd9))))?((-4'sd0)?(4'sd3):(-2'sd0)):((5'd21)?(5'sd9):(4'sd4))))));
  localparam signed [3:0] p3 = (((2'sd0)?(5'sd6):(2'd3))?((5'sd15)?(-4'sd4):(2'd2)):((2'd0)?(3'd3):(5'd19)));
  localparam signed [4:0] p4 = ((((2'd2)>(5'd17))<=((3'd1)?(2'sd0):(5'd1)))&((~|((2'sd0)?(2'd2):(3'd6)))==={4{(-3'sd3)}}));
  localparam signed [5:0] p5 = (({(2'd1),(2'sd1),(3'd1)}>>{(4'd15)})&((~&(-3'sd0))-((2'd0)^~(-2'sd0))));
  localparam [3:0] p6 = ((-4'sd1)>=(-4'sd1));
  localparam [4:0] p7 = {((+(((-4'sd0)>>>(-4'sd2))|((4'd15)+(4'd4))))<(+((&(-4'sd5))&&(~&(5'd20)))))};
  localparam [5:0] p8 = (2'sd1);
  localparam signed [3:0] p9 = ((((2'sd0)^(-5'sd7))!=((5'sd8)?(5'd19):(5'sd5)))&&(((4'd14)/(5'd27))>>(|((2'd1)&&(4'sd0)))));
  localparam signed [4:0] p10 = {3{{1{{1{{1{(3'd6)}}}}}}}};
  localparam signed [5:0] p11 = ((~^((^(~&(2'd0)))-((2'sd0)^~(-4'sd6))))^~(+((~&((5'd13)===(5'sd5)))!==(~&((-2'sd1)<(4'sd3))))));
  localparam [3:0] p12 = ((~|(&(~&{(-4'sd2),(4'sd0),(2'd0)})))-{((-3'sd1)^(2'sd1)),{4{(3'd3)}}});
  localparam [4:0] p13 = ((&((2'd0)===(2'sd1)))-((-4'sd0)?(4'sd5):(4'd5)));
  localparam [5:0] p14 = (((-5'sd9)&(-3'sd3))>=((-3'sd2)>>(-4'sd2)));
  localparam signed [3:0] p15 = (~((6'd2 * {2{(3'd4)}})<((3'sd3)>={3{(2'd0)}})));
  localparam signed [4:0] p16 = (4'd13);
  localparam signed [5:0] p17 = {(~^(3'd1)),(+(4'd6)),(3'sd3)};

  assign y0 = (&(|$unsigned(((b0===b5)^~$unsigned(p11)))));
  assign y1 = ((-(~^(-4'sd7)))-($unsigned((~|b1))?(b5?p5:p2):(a1-a1)));
  assign y2 = (~&(-5'sd12));
  assign y3 = {1{({3{(p7?a3:p17)}}?{4{p0}}:((p16?p0:p16)?(5'sd10):(p3?p10:p4)))}};
  assign y4 = (4'd15);
  assign y5 = {(~&{(p1?b0:a3)}),(^(!$signed(a4)))};
  assign y6 = (4'd3);
  assign y7 = (({3{a5}}|(b3&b5))&{1{((a1<a4)!==(b5>=b1))}});
  assign y8 = {{{(~&{4{b2}})}},{4{(&a5)}}};
  assign y9 = {3{(a0||p2)}};
  assign y10 = (((p14<<<p17)>=(6'd2 * a2))>=((b2||b5)!=(a3>=b4)));
  assign y11 = ((^($signed(b5)?(~&a0):(a5)))?((a0)?(|b4):$unsigned(a4)):($signed(p9)?(b1?b2:a1):(a2?p2:b5)));
  assign y12 = (5'd2 * (!(p6<<<p8)));
  assign y13 = (({4{b4}}-(~b2))?(~(a3<=a4)):(a2?a5:b4));
  assign y14 = (~&(4'd7));
  assign y15 = ({{a5,p7,p11},{b0},(-4'sd3)}+(4'd8));
  assign y16 = ((a3>=b1)?{2{p16}}:{4{a5}});
  assign y17 = ((-2'sd1)&&(~(p17?p9:p3)));
endmodule
