module expression_00697(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (({(-5'sd2)}!=={3{(-4'sd1)}})>>>(~|{{4{(-4'sd2)}}}));
  localparam [4:0] p1 = (((-4'sd0)/(-5'sd7))<=((-4'sd6)===(-4'sd3)));
  localparam [5:0] p2 = (((~|(~^{2{(-5'sd5)}}))<((4'd12)^((-4'sd5)!==(-5'sd12))))&&(5'd1));
  localparam signed [3:0] p3 = (((3'd4)?(-5'sd11):(5'sd3))?(((-3'sd0)|(4'd4))<((-5'sd6)>(5'd28))):(4'd6));
  localparam signed [4:0] p4 = ((!(-(~((4'sd4)>>>(4'sd3)))))?(((5'd28)?(4'd12):(5'd10))?{4{(3'd7)}}:{4{(-4'sd0)}}):{3{{4{(4'd14)}}}});
  localparam signed [5:0] p5 = ((((4'sd6)<(5'sd11))=={(-4'sd2),(3'd2)})<<<{{2{(4'd6)}},{(2'd1)},(2'sd0)});
  localparam [3:0] p6 = (-3'sd2);
  localparam [4:0] p7 = {(2'sd0),(|((-4'sd4)-(3'sd3)))};
  localparam [5:0] p8 = (5'd24);
  localparam signed [3:0] p9 = (~|({((4'd14)!==(5'd7)),(!(4'd8)),(~&(4'd11))}||((~|((5'sd0)+(4'd3)))^~(2'd1))));
  localparam signed [4:0] p10 = ((~^(6'd2 * ((2'd3)<<<(2'd1))))>=((^(&(4'sd0)))>(~((4'sd2)?(-5'sd10):(2'sd0)))));
  localparam signed [5:0] p11 = (4'd6);
  localparam [3:0] p12 = {(~&(2'd1)),((2'd2)<<<(-3'sd1)),(4'sd2)};
  localparam [4:0] p13 = (^(~|(&{(^((+(4'd6))===(~^(-3'sd2)))),(&(~(~(-(2'sd1)))))})));
  localparam [5:0] p14 = (2'sd1);
  localparam signed [3:0] p15 = {3{((-5'sd3)|{1{(3'd0)}})}};
  localparam signed [4:0] p16 = ({(-4'sd6),((-4'sd5)>=(2'd2)),((2'd0)<(2'd1))}?(-3'sd2):{(3'd4),(3'sd2),((5'sd13)?(4'd5):(2'sd0))});
  localparam signed [5:0] p17 = {2{(2'd2)}};

  assign y0 = (~|(!((~(b2<<<a3))*(b5===a3))));
  assign y1 = (2'd0);
  assign y2 = {1{(~&p10)}};
  assign y3 = (^((^{(~^((-b1)!=(~^a2)))})|((|(~|$signed(a5)))<({p14,b4,a4}>>>(+a4)))));
  assign y4 = {2{(p12||b4)}};
  assign y5 = ((((b2!=a1)))<<((3'sd1)==={3{b5}}));
  assign y6 = (!{2{(-{a1,a4,a4})}});
  assign y7 = ((b3>>>a0)!=(+a2));
  assign y8 = {4{{{2{b3}},{2{a3}}}}};
  assign y9 = (^((~&(b1?p12:b1))==(p11?p3:p17)));
  assign y10 = {4{$unsigned((b0>>>p10))}};
  assign y11 = ((b3+a5)===(a2^~b3));
  assign y12 = {((p0==p10)&&{p0}),((a2==b5)===(b0>b2))};
  assign y13 = ({p3,b5}?(p17^~p9):(~^a2));
  assign y14 = ({2{(p12?p10:b5)}}?$signed((p8?p3:p4)):((b2&&p11)-$signed(p17)));
  assign y15 = {((4'sd0)&&(2'd0))};
  assign y16 = (~|({(b1<<p10),(~p17),(p4>=p17)}>($signed(b4)^(p2>p1))));
  assign y17 = (+(~^(!(^(-(^(~(~&(!(~(~(|(~|(|(~|(~&p2))))))))))))))));
endmodule
