module expression_00635(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (3'd2);
  localparam [4:0] p1 = ((^((4'd15)<(-5'sd5)))+{(~(-4'sd4)),{4{(-2'sd0)}}});
  localparam [5:0] p2 = ((3'sd1)?(3'd5):(-5'sd1));
  localparam signed [3:0] p3 = ((|{3{(2'd3)}})?((~(-4'sd6))?{3{(2'd3)}}:{2{(4'd3)}}):(((4'd4)?(5'd19):(5'd3))?((3'd5)>=(4'sd7)):{4{(5'sd2)}}));
  localparam signed [4:0] p4 = (-(-4'sd2));
  localparam signed [5:0] p5 = ((6'd2 * ((4'd8)>=(4'd12)))<<({(4'd2)}&&((2'd2)<<(2'd0))));
  localparam [3:0] p6 = (~&(3'sd0));
  localparam [4:0] p7 = (2'd2);
  localparam [5:0] p8 = ((~|(5'sd8))<<(4'd12));
  localparam signed [3:0] p9 = (-((5'd27)^(4'sd2)));
  localparam signed [4:0] p10 = ((-{4{(2'sd0)}})>>>((4'd9)>>>(2'd3)));
  localparam signed [5:0] p11 = {((4'd14)?(3'd1):(3'd3)),((4'd8)?(-5'sd3):(5'sd3)),((5'sd4)+(4'd1))};
  localparam [3:0] p12 = {4{((2'sd0)^~(-3'sd2))}};
  localparam [4:0] p13 = (((-2'sd0)<=((-4'sd4)-(3'sd1)))&(((-3'sd2)>=(3'd0))>>(~^(-3'sd2))));
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = ((2'd1)?(3'd7):(-5'sd7));
  localparam signed [4:0] p16 = ((~|{4{(3'd5)}})&&(4'sd7));
  localparam signed [5:0] p17 = (6'd2 * (2'd0));

  assign y0 = (p3!=a3);
  assign y1 = (-(&{(a5>=b1),(-a5),(b5!=b0)}));
  assign y2 = ((5'sd9)>(~((4'sd5)>>(2'd2))));
  assign y3 = (2'd3);
  assign y4 = (&(((p12&p3)?(a1>>a4):{a3,a0,a0})&&(~|(+((a0==b2)&&(~b2))))));
  assign y5 = (((5'd2 * p0)-(4'd2 * b1))||((b3<=a0)-(p4!=a4)));
  assign y6 = (-3'sd1);
  assign y7 = (^(+{3{p17}}));
  assign y8 = (((((b3<=a2)))===$unsigned((a1^~b3)))||($signed(($signed(((p5<<p5)>(a0>p15)))))));
  assign y9 = {(({b2}<(p0^~p5))>=({4{p6}}<<{1{p2}})),{((b4&a5)==={3{b1}}),{2{(p4)}}}};
  assign y10 = (!{a3,a2,a1});
  assign y11 = (({({p16,p11}>=(p9-p2))}>=((p17&&p17)>>>(^p13)))<<(((~p12)>=(2'd1))<(~^((p14<<<p4)>(p10<<<p8)))));
  assign y12 = {2{(b3!=b5)}};
  assign y13 = {3{(-3'sd1)}};
  assign y14 = (((b1?a4:a0)||(b5?b3:b5))?((a0?b5:a3)?(6'd2 * a0):(b5&b1)):((b2>=b5)|(6'd2 * b0)));
  assign y15 = (2'd2);
  assign y16 = {2{(3'sd1)}};
  assign y17 = $unsigned({{1{{$signed({{1{{2{{{3{b1}},{4{b5}},{1{b5}}}}}}}})}}}});
endmodule
