module expression_00883(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'd3)>=(-2'sd0))*((2'd2)-(-4'sd7)))!==(((5'd17)===(4'sd0))===((-2'sd1)!==(3'd4))));
  localparam [4:0] p1 = (6'd2 * ((3'd1)&(2'd2)));
  localparam [5:0] p2 = (!{2{(5'd27)}});
  localparam signed [3:0] p3 = (^{(~^(5'd26)),{2{(-2'sd1)}},((2'sd1)==(-5'sd4))});
  localparam signed [4:0] p4 = ({{(5'd26),(5'd30),(5'sd10)},{2{(-2'sd0)}}}?(~^((4'd15)?(2'd3):(5'sd14))):(!(^{4{(3'd1)}})));
  localparam signed [5:0] p5 = {{(+(4'sd4)),(~(-2'sd1))},{4{(-2'sd0)}},{3{{3{(2'd1)}}}}};
  localparam [3:0] p6 = (((4'd12)>>>(4'sd5))/(-5'sd13));
  localparam [4:0] p7 = ((((5'd0)||(-4'sd5))<<(4'sd1))>>>(((5'd24)?(-4'sd2):(4'd5))===((-2'sd1)?(2'd3):(5'd31))));
  localparam [5:0] p8 = (((2'd1)||(5'sd7))+((2'd2)*(2'd3)));
  localparam signed [3:0] p9 = ({3{(4'd0)}}|(3'sd2));
  localparam signed [4:0] p10 = (^((+((3'd4)?(5'd16):(2'd3)))?((2'sd0)?(-5'sd13):(5'd7)):((5'sd0)?(-3'sd0):(4'sd2))));
  localparam signed [5:0] p11 = ({4{(2'd0)}}>>(((5'd17)|(-4'sd5))==(4'd8)));
  localparam [3:0] p12 = ((^(&(~&(((3'd1)&(2'sd1))<<<(-(5'sd13))))))&&(((3'sd3)^(2'd2))<<<((5'sd0)!==(2'd3))));
  localparam [4:0] p13 = {2{{1{((5'sd0)?(4'sd7):(-4'sd2))}}}};
  localparam [5:0] p14 = ({2{(2'd1)}}&((3'd2)>>(2'd2)));
  localparam signed [3:0] p15 = ((5'd25)<=(4'd6));
  localparam signed [4:0] p16 = (!{2{(4'd8)}});
  localparam signed [5:0] p17 = {(!(2'd0)),(+(4'd13))};

  assign y0 = (~&((-(~^{(~|p6),{b3,a4,p1},(~|p6)}))-(|{((~|(!a0))!={p15,b0,p2})})));
  assign y1 = (!(~&(-(~(((!{a5})!=$unsigned((|b0)))>>$unsigned({(a3^b0),(+b4),{b2}}))))));
  assign y2 = (!((!(p11^~a5))>=((p16|p10)<<<(-b1))));
  assign y3 = (-{2{{4{b3}}}});
  assign y4 = {3{$signed(({4{a4}}==(p2)))}};
  assign y5 = (5'd16);
  assign y6 = (|{3{(~(-5'sd4))}});
  assign y7 = (4'd2 * (p1?p7:p12));
  assign y8 = (^(!{(~|((!((|b4)?(~^p9):(a3?a2:p14)))?(|({a2,a0}?(&b4):(^b5))):(~&((a3?b3:p0)?(p9?a1:b4):(~a4)))))}));
  assign y9 = {(($signed(p9))!=(b0!==a5)),(-(~(3'd6)))};
  assign y10 = ({(&(|({1{(b0!==a2)}}<<<(~{3{b0}}))))}^~(&(((b5?b4:a0)!=(a5<<a4))==={3{b2}})));
  assign y11 = (~&{(~{(~&(-p13)),{p8,b0}}),(~^(|(~^{{p17,p12},(~^p1)})))});
  assign y12 = (-5'sd11);
  assign y13 = {{((3'd0)?(5'sd14):{3{a3}})},((a4&&b0)?(5'sd3):(b3?a4:a4))};
  assign y14 = {3{{3{p12}}}};
  assign y15 = (|(~|(a4||a3)));
  assign y16 = ((-((+(3'd5))%a5))<<<(-(~&(|((~p6)&&(~^p5))))));
  assign y17 = (-{(!(^(~{((!(-a5))<<<$unsigned((&p4)))})))});
endmodule
