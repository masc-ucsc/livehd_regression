module expression_00733(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd1)?(5'd25):(-5'sd3))?(~((5'd13)?(5'd7):(5'd10))):(-2'sd1));
  localparam [4:0] p1 = ((4'd6)?(4'd1):(-2'sd0));
  localparam [5:0] p2 = (((3'sd0)?(-2'sd0):(4'd2))?((5'sd11)?(-5'sd12):(-3'sd2)):(~^(4'sd0)));
  localparam signed [3:0] p3 = (~{((3'd1)?(2'd3):(2'd3)),(5'd2 * (4'd7)),((2'sd1)===(4'd8))});
  localparam signed [4:0] p4 = ({3{(-5'sd7)}}<<{1{((3'sd3)>(5'd31))}});
  localparam signed [5:0] p5 = {(((5'sd0)?(-5'sd13):(3'sd2))?(^((4'sd5)?(2'd1):(3'd5))):((3'd0)?(3'sd0):(-4'sd5)))};
  localparam [3:0] p6 = ((-((-2'sd0)?(3'sd0):(-5'sd2)))&&(!((3'd7)||((3'd7)^(2'd1)))));
  localparam [4:0] p7 = {{(({(3'sd2)}?{(3'd7)}:((-5'sd14)?(3'd4):(-5'sd2)))===(((-2'sd0)==(2'd0))>={(&(3'sd3))}))}};
  localparam [5:0] p8 = (5'd2 * {1{(~(4'd3))}});
  localparam signed [3:0] p9 = (~|({(-4'sd6),(-2'sd1),(-2'sd0)}|{(-2'sd0),(2'd2)}));
  localparam signed [4:0] p10 = {({((3'sd0)?(2'd1):(5'd11)),{(4'd5),(2'd3),(5'sd1)},{(4'sd3),(4'd3),(-2'sd0)}}?{((-5'sd14)?(2'd1):(-5'sd2)),((4'd13)?(5'd16):(3'd0)),{(2'd2)}}:(((4'sd4)?(2'sd1):(3'd5))?((-5'sd0)?(2'sd0):(5'sd3)):((2'sd0)?(3'd5):(3'd4))))};
  localparam signed [5:0] p11 = ((-3'sd3)<=(3'd6));
  localparam [3:0] p12 = (~|({1{{1{(3'd5)}}}}>=(+((3'd6)>>>(5'sd8)))));
  localparam [4:0] p13 = (4'sd3);
  localparam [5:0] p14 = (((-5'sd13)>(-3'sd0))<<((4'sd7)===(5'd17)));
  localparam signed [3:0] p15 = {{(5'sd0),(3'd1),(-4'sd0)},{{(3'sd0),(4'd2),(-4'sd5)},{(3'd1),(-4'sd1)}},(~^(~|(~&(-5'sd1))))};
  localparam signed [4:0] p16 = (~&(((2'd1)/(-5'sd1))|(5'd6)));
  localparam signed [5:0] p17 = (~{((~&(4'sd6))?(~(2'sd1)):(~(3'd5)))});

  assign y0 = ((({4{b2}}<=(!p14))>{3{(b5?b1:b3)}})>>(((p6|p0)?(~^a0):{3{a0}})<({a1,p4,a2}||{b3,a5})));
  assign y1 = (^{(2'sd0)});
  assign y2 = {((a3<<<b5)+(b1>a0)),(5'd2 * {b2,a2}),((b1<a4)<{b2,a5})};
  assign y3 = ((~^(4'd5))?(~^((p6>p8)|(|p6))):((p10?p16:p9)?(b1+p16):(p11?p12:p13)));
  assign y4 = {2{b5}};
  assign y5 = ((~|(p14?a0:a3))<<<((b4|b3)*(~&b4)));
  assign y6 = (|(((b4)?(b2?b5:b0):{2{p4}})?($unsigned(b3)?(b2==a3):(+a2)):((b1>=a2)?$signed(p14):{3{b4}})));
  assign y7 = {2{$signed((~&(p4<=a2)))}};
  assign y8 = {2{{4{a2}}}};
  assign y9 = {1{(({b1,b5}&&{4{b4}})&&(!((~&{a5,a1})+(a4>=a1))))}};
  assign y10 = $signed((5'd17));
  assign y11 = (5'd2 * (a0<<a2));
  assign y12 = (+((((^b3)>=(p11-b3))>>((a1+a4)+(b0)))|(((b2|p10)^~(p4))-((a4&&b0)))));
  assign y13 = {(a4>>p14)};
  assign y14 = (!(+(~^((-a4)?{p5}:(|a1)))));
  assign y15 = ((p14>>p8)-(5'd25));
  assign y16 = {1{((p9<<a2)?(a1>=a3):(b5?b5:a4))}};
  assign y17 = (a0<p0);
endmodule
