module expression_00943(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'd2)?(2'd2):(-5'sd5))&&((3'd2)?(-2'sd0):(2'd3)))+(((3'd6)?(4'sd2):(3'd1))<=((3'd2)?(2'sd1):(3'd7))));
  localparam [4:0] p1 = (2'sd0);
  localparam [5:0] p2 = (~^((|{(5'sd10),(5'sd9)})?(-{(-4'sd6),(5'sd10),(4'd14)}):(~&((3'd4)?(2'd3):(2'd0)))));
  localparam signed [3:0] p3 = (&{(((3'd0)>=(4'd3))+{(4'd15),(3'd6)}),{((5'sd8)&&(2'd0))},{(-(2'd2)),((2'sd0)<=(-2'sd0))}});
  localparam signed [4:0] p4 = ((4'd10)===(2'd1));
  localparam signed [5:0] p5 = (((-2'sd0)?(3'd7):(3'd5))?{2{(4'd7)}}:((3'd0)<<(3'sd2)));
  localparam [3:0] p6 = (3'sd3);
  localparam [4:0] p7 = {3{(&(~&(-((-2'sd1)&(5'd21)))))}};
  localparam [5:0] p8 = (-3'sd2);
  localparam signed [3:0] p9 = ({{4{((-4'sd4)!==(-5'sd5))}}}+(((-3'sd1)?(5'sd3):(5'sd14))>(((3'd6)<=(5'd31))>={(3'd4),(5'sd7)})));
  localparam signed [4:0] p10 = (&(5'sd0));
  localparam signed [5:0] p11 = (~^(({3{(-2'sd0)}}+((3'd6)?(3'd7):(3'd4)))?(((5'sd8)==(2'd0))?((5'd19)<<<(4'sd2)):((2'd1)?(2'sd0):(-5'sd7))):((2'd2)>>>{2{(3'd1)}})));
  localparam [3:0] p12 = {(!(+{(4'sd4),(-2'sd0),(5'sd1)})),{4{(2'd3)}},(~|(3'd4))};
  localparam [4:0] p13 = {3{{2{(2'sd0)}}}};
  localparam [5:0] p14 = {3{{1{(5'd22)}}}};
  localparam signed [3:0] p15 = (((3'd3)>>(-5'sd8))?((3'd5)!=(4'sd1)):((-3'sd0)<=(4'd13)));
  localparam signed [4:0] p16 = (6'd2 * (5'd31));
  localparam signed [5:0] p17 = {(!{{(-2'sd0),(3'd1),(5'd7)},{(2'd0),(3'd5)},((-3'sd3)!=(3'd2))})};

  assign y0 = (+(((2'd0)>{1{b5}})<=((2'd1)!=(b2?b4:p13))));
  assign y1 = (^{2{(3'sd3)}});
  assign y2 = (({{4{a5}}}^((a3<<<p3)^~(a3|b3)))<((b5?p13:p13)?({p17}):$unsigned((a3<<<b0))));
  assign y3 = (5'd2 * (b1===b1));
  assign y4 = $signed({(|{p10,p2,p15}),(!$signed((-p14)))});
  assign y5 = {4{p13}};
  assign y6 = ((~&(|((p5?a1:a4)&&(~a5))))?(-{4{b1}}):{1{{1{(p7?a4:a3)}}}});
  assign y7 = (3'd7);
  assign y8 = (a1<<a2);
  assign y9 = {2{b0}};
  assign y10 = {((a1!==b1)>=(b3&b4))};
  assign y11 = ((-5'sd5)+{(a0?a1:a1),(4'd2 * a2)});
  assign y12 = (2'd0);
  assign y13 = {(5'sd8)};
  assign y14 = (a1?a1:p10);
  assign y15 = (~^(p1?b1:a1));
  assign y16 = (&(4'd2 * (|(b1*b2))));
  assign y17 = ((^({1{(~p5)}}<<{p4,p5,p10}))<<(-({1{(b4!==a5)}}>=(p6!=p6))));
endmodule
