module expression_00130(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^(~(&(3'd1))));
  localparam [4:0] p1 = (|{(~&(|(~^(~|{(-(5'd5)),((3'd2)>(2'sd0)),(|(4'd2))}))))});
  localparam [5:0] p2 = ((((3'sd0)>>>(2'd2))||((4'd9)>>>(4'sd6)))<<(5'd2 * (~((3'd5)?(2'd2):(4'd12)))));
  localparam signed [3:0] p3 = (5'd21);
  localparam signed [4:0] p4 = (~&{(~^(-3'sd3))});
  localparam signed [5:0] p5 = (&(^(+(~^(&(~|(+(^{{(5'sd13),(-3'sd2),(2'd0)},(|(3'd4))}))))))));
  localparam [3:0] p6 = (~&(3'd5));
  localparam [4:0] p7 = (4'd4);
  localparam [5:0] p8 = {2{(~^{(2'd2),(4'd1)})}};
  localparam signed [3:0] p9 = {(!((-5'sd2)>(4'd0))),{((-2'sd1)===(4'd9)),((2'd3)<<<(3'sd0))},(+(^((-3'sd2)<<<(5'd11))))};
  localparam signed [4:0] p10 = (|((3'sd2)?(4'd15):(5'sd13)));
  localparam signed [5:0] p11 = {1{({2{(4'sd4)}}|((5'sd11)>>(4'd11)))}};
  localparam [3:0] p12 = (((3'd6)==(2'd3))||(!(-(3'sd2))));
  localparam [4:0] p13 = ({(4'd7),(2'd0),(2'd1)}<=((-2'sd1)||(2'd3)));
  localparam [5:0] p14 = ((((-2'sd0)?(3'sd3):(-2'sd1))?(|(4'sd7)):{1{(3'd2)}})^~((~^(2'sd1))?((5'd9)^~(-4'sd7)):(|(-5'sd11))));
  localparam signed [3:0] p15 = {2{(5'sd15)}};
  localparam signed [4:0] p16 = (-{((5'd18)>=(-2'sd0))});
  localparam signed [5:0] p17 = ({{(3'd6),{4{(4'd12)}}},({1{(5'd29)}}^(!(3'd4)))}||(~|({(-4'sd6),(5'd20),(2'd0)}>=((2'sd1)|(-2'sd1)))));

  assign y0 = (5'd2 * (a0<=a0));
  assign y1 = (p4?a2:b3);
  assign y2 = {(~(-2'sd1))};
  assign y3 = (&(&a3));
  assign y4 = {4{{1{p13}}}};
  assign y5 = ((b4?a2:a0)!==(a0?b1:b4));
  assign y6 = ($signed(({$unsigned(p1),{a1,p1,a4}}&&({a3}||(a1>p16))))==($signed({$unsigned({b1,a4})})==={((a0>>b2)>>>(b1<=a0))}));
  assign y7 = $signed(((2'd0)));
  assign y8 = {(!(({a2,b1,b2}===(~&(~(b2<=b1))))&&(({a0,a3}&(&p6))<{(b4!==b2),(~^b3)})))};
  assign y9 = (-2'sd1);
  assign y10 = (((-a4)|(~&b1))===({1{b2}}>={1{b5}}));
  assign y11 = {$unsigned($signed($unsigned(p1))),{($unsigned(p13))}};
  assign y12 = (&((p12+p2)>(~|{p6})));
  assign y13 = ((a5===a3)>=(4'sd1));
  assign y14 = $unsigned((~|$signed(b5)));
  assign y15 = (((+b5)?(-a2):(-p9))?(6'd2 * (p2+p1)):((p8%b0)?(~|p7):(p11/p11)));
  assign y16 = (-(2'sd1));
  assign y17 = ((-2'sd0)==({2{{1{p3}}}}^~(2'd3)));
endmodule
