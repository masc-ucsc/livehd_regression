module expression_00048(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (^(4'sd1));
  localparam [4:0] p1 = ({((3'd7)?(5'sd12):(2'd3)),{1{(-2'sd1)}}}?{{(-2'sd1)},((3'sd1)==(2'd0))}:{4{(3'd5)}});
  localparam [5:0] p2 = ({(2'd2),(4'd7)}&&((4'd10)>>(4'd8)));
  localparam signed [3:0] p3 = (((4'd8)!==(4'd0))|((3'd6)||(-3'sd2)));
  localparam signed [4:0] p4 = ((2'd1)?(4'd8):(2'sd1));
  localparam signed [5:0] p5 = {2{(3'd3)}};
  localparam [3:0] p6 = (((2'd1)-((-5'sd10)!=(5'sd13)))<=(-(|(~((4'd10)<<<(3'sd1))))));
  localparam [4:0] p7 = ((5'd2 * ((4'd8)^(3'd7)))!=({(5'sd11),(4'd11),(4'sd6)}<=(~^(3'd6))));
  localparam [5:0] p8 = (~|(+((+(4'd2 * (2'd1)))|((5'd14)<(2'd2)))));
  localparam signed [3:0] p9 = (((-3'sd0)?(2'sd0):(4'd1))^(~^(-3'sd0)));
  localparam signed [4:0] p10 = ((-3'sd2)?(2'd2):(5'd22));
  localparam signed [5:0] p11 = (4'd13);
  localparam [3:0] p12 = {3{{4{(2'd3)}}}};
  localparam [4:0] p13 = (!{{(5'd29),(3'd3)},{3{(5'd20)}}});
  localparam [5:0] p14 = (((4'd7)===(2'sd1))*((5'd3)?(5'd29):(2'd1)));
  localparam signed [3:0] p15 = ((-4'sd5)?(4'd7):(((4'd7)?(3'd1):(-4'sd0))<<<((4'sd1)>(4'd5))));
  localparam signed [4:0] p16 = ((2'sd0)&&(3'sd2));
  localparam signed [5:0] p17 = ((2'd1)-(3'd6));

  assign y0 = $unsigned(((~&(~&(4'd2 * p12)))));
  assign y1 = (3'd1);
  assign y2 = $signed({4{{1{((b0^a4))}}}});
  assign y3 = (!($signed(a0)?$signed(b0):(p5>>>p0)));
  assign y4 = (6'd2 * $unsigned((p10>>p6)));
  assign y5 = (~|({3{(~^p17)}}^{{4{p15}},(~&p16),(b3!==b2)}));
  assign y6 = (!{1{$signed(({3{$unsigned((&{4{p15}}))}}))}});
  assign y7 = (|(~$signed(((-5'sd1)-{4{b5}}))));
  assign y8 = (-4'sd1);
  assign y9 = (-(+(~|{$signed({({(|b0),(5'sd6)}),(3'sd3),(5'sd10)})})));
  assign y10 = $unsigned($signed((4'd15)));
  assign y11 = (b0<a4);
  assign y12 = ((^(~&(~|(-5'sd5))))>=((-p5)>(b1!==a2)));
  assign y13 = ($unsigned(((p1<<<p15)||(p17)))?((a1?b3:p8)?(p4):(p8&p6)):$unsigned(((p16?p12:p4)^~(4'd2 * a0))));
  assign y14 = {a0,p5,p1};
  assign y15 = {4{{(+a5),{4{p6}},(b3>>>a5)}}};
  assign y16 = (~&{({p3,p2}==(a1&p13))});
  assign y17 = ((~&(b0<<<a5))>(b2-b5));
endmodule
