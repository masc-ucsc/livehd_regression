module expression_00553(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ({4{(4'd6)}}-((+(-2'sd0))<<{3{(3'sd1)}}));
  localparam [4:0] p1 = (((|(~^(2'd2)))||((-5'sd12)^(3'd7)))!=((~|(^(5'd1)))<<((5'sd11)<=(-5'sd8))));
  localparam [5:0] p2 = (3'sd1);
  localparam signed [3:0] p3 = (((3'sd0)?(5'sd3):(4'd4))?{4{(-4'sd6)}}:{3{(-5'sd10)}});
  localparam signed [4:0] p4 = ((((4'd3)^~(2'd3))^~((3'd0)==(5'd7)))?(((-2'sd1)?(3'd3):(3'd7))>((-2'sd0)<(5'sd6))):((-5'sd3)?(4'sd4):(4'd8)));
  localparam signed [5:0] p5 = (3'd6);
  localparam [3:0] p6 = ({(-5'sd4),(-3'sd0)}-(!(2'd1)));
  localparam [4:0] p7 = {{(2'd1),(2'd1),(5'd20)},{4{(2'd3)}}};
  localparam [5:0] p8 = (({(-2'sd0),(4'd12),(-4'sd4)}>>>((5'sd13)||(5'd31)))==(4'd2 * {2{(5'd18)}}));
  localparam signed [3:0] p9 = {(2'sd1),(3'd3),(5'sd0)};
  localparam signed [4:0] p10 = (2'd1);
  localparam signed [5:0] p11 = ((+(-(4'd5)))>=((5'd2)?(2'd0):(4'sd1)));
  localparam [3:0] p12 = ((~^(~(~^((2'd2)?(4'sd1):(-5'sd4)))))<<((~|(2'sd1))?((4'sd7)?(4'd7):(2'sd1)):((-5'sd5)^~(-3'sd1))));
  localparam [4:0] p13 = (((3'd1)!==(-4'sd0))*((-4'sd4)&(2'sd1)));
  localparam [5:0] p14 = (~^(((+(~^(-3'sd2)))!=((4'd0)>(2'd3)))&&{((4'd0)>=(3'sd0)),(4'sd6)}));
  localparam signed [3:0] p15 = ((3'sd3)||(3'd6));
  localparam signed [4:0] p16 = (~^((-2'sd1)!=(-2'sd0)));
  localparam signed [5:0] p17 = {(4'd15)};

  assign y0 = ($signed({1{((~|p2)-$unsigned(a5))}})<<<({1{(~&b3)}}<(&(^a4))));
  assign y1 = $signed({1{(({3{(a1)}})!==({4{b3}}^~({a0})))}});
  assign y2 = (((a3?a1:b4)==(a2<p13))^~(-(a2?b0:b4)));
  assign y3 = (5'd2 * {p2,p7,p6});
  assign y4 = ((-5'sd9)!==({3{b1}}&&(b5>=a4)));
  assign y5 = (!(((({p6,a0,a4}<<(p9^a0))-{(p1==p1)}))));
  assign y6 = (a3?a0:b0);
  assign y7 = ((-5'sd15)+{4{p9}});
  assign y8 = {((b2?p7:p8)?(2'd0):{b2}),((a3?p15:a1)?(p4>>a1):{p9}),((~|p15)&(-4'sd1))};
  assign y9 = ((b4<<b2)!=(~(2'd2)));
  assign y10 = {3{(p10<<p12)}};
  assign y11 = (p3?p11:p11);
  assign y12 = $signed({4{{1{{$signed(a0),{1{b4}}}}}}});
  assign y13 = {3{p7}};
  assign y14 = (((-5'sd1)+((a2>>b3)===(~^a3)))^(3'd0));
  assign y15 = $unsigned({(a3?p7:p0)});
  assign y16 = {1{((&{2{{{a3,a5}}}})-((|(a0>>>b0))>((~&(!b4)))))}};
  assign y17 = (b1&b0);
endmodule
