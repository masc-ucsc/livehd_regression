module expression_00864(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(~((|(|(4'd7)))&((-(5'd31))^((-4'sd1)!=(-5'sd1))))));
  localparam [4:0] p1 = ({(3'sd0)}?{{(5'sd1),(5'sd0),(3'd6)}}:{(5'd4),(2'd0)});
  localparam [5:0] p2 = (((-3'sd2)<<<(5'd17))<=(!((5'd17)*(4'sd3))));
  localparam signed [3:0] p3 = (((4'sd0)<<(-3'sd2))<<((2'd3)&(4'd13)));
  localparam signed [4:0] p4 = ((|(4'sd4))?(&(5'sd10)):{(3'd6),(4'd11)});
  localparam signed [5:0] p5 = (3'd7);
  localparam [3:0] p6 = {((&(5'sd1))|((5'd29)<(3'd6))),(~|(~{(3'd1),(3'd3),(5'd18)}))};
  localparam [4:0] p7 = ((2'd2)&{((-2'sd1)|(4'd2)),(4'd2 * (5'd9))});
  localparam [5:0] p8 = (2'd2);
  localparam signed [3:0] p9 = (((3'sd3)+(-5'sd0))?((3'd0)&(4'sd2)):((4'd14)?(5'sd1):(2'd2)));
  localparam signed [4:0] p10 = ((((-3'sd0)%(3'sd3))>=((4'd7)%(-3'sd0)))-(((-2'sd0)==(-4'sd2))!==((5'd4)!=(2'd0))));
  localparam signed [5:0] p11 = (~((&(((5'd9)<=(5'd23))||(-(4'd11))))^(((4'd3)>>>(3'd0))||((2'd3)^~(3'sd3)))));
  localparam [3:0] p12 = (~|(!(((2'd3)?(2'd0):(-3'sd3))?(~((5'sd0)?(-4'sd2):(3'sd2))):((-5'sd1)?(2'd1):(-4'sd5)))));
  localparam [4:0] p13 = ((~^((-2'sd1)>=(4'sd7)))!=(-((-3'sd2)<<(-5'sd5))));
  localparam [5:0] p14 = (&(!(4'sd1)));
  localparam signed [3:0] p15 = (((2'sd0)^~(4'sd5))>{(2'd3),(5'd21),(5'd12)});
  localparam signed [4:0] p16 = (({1{{(-2'sd1),(2'd0),(4'd4)}}}^~{(3'd2),(3'd7)})>({(2'd3),(2'd0)}^~{(2'd3),(4'd7),(3'sd2)}));
  localparam signed [5:0] p17 = ((2'd0)!==(4'd6));

  assign y0 = (({2{(~|a4)}}>>{{p3,p5,a0},{3{p0}}})&&(^(((~|p13)>={1{p2}})^((b5+a1)>=(p8&&p9)))));
  assign y1 = {(2'd3),{($signed(b2)),(&(p3))},{(^{a4,p9,b1})}};
  assign y2 = (+(b3*p11));
  assign y3 = {((p4>=p4)&&(p2^p11)),{(p13<=p9)},((5'sd7)>=(p6))};
  assign y4 = ((p10?p8:a2)?{1{{2{p2}}}}:(&(4'd11)));
  assign y5 = (p2>>>p1);
  assign y6 = ((((-2'sd1)>(6'd2 * b0))<={2{(3'sd2)}})&&(+((b0||b2)!=(!(b1!=a3)))));
  assign y7 = ({(p16?b4:b3),(~|{1{b3}})}==((!(~a2))<={p7,p8,a1}));
  assign y8 = {{{p0},{p0,a3,p12},{p11}},{(a3?p3:a5),{(a1?p17:a4)}},{(a5?p8:p14),{p14,a1,p8}}};
  assign y9 = ({p14,p4}?((3'd1)):((p10?p6:p5)));
  assign y10 = (2'd1);
  assign y11 = {1{a5}};
  assign y12 = {{2{a0}},{2{b2}}};
  assign y13 = {2{(2'd3)}};
  assign y14 = (|(!($unsigned(a3)?$signed(a5):$unsigned(b0))));
  assign y15 = (4'd1);
  assign y16 = (|(~((((2'd1)&&$signed((p9<<p6)))>>>((-(a5?b3:b1))!==(b1?a4:b4))))));
  assign y17 = {(((b5!==b0)-{(b3+b0)})!=={{b4,b2,b2},{a3,b5,b2},(b4>b2)})};
endmodule
