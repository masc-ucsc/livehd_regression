module expression_00541(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-4'sd1);
  localparam [4:0] p1 = ({1{(^{2{{4{(-4'sd7)}}}})}}^~({2{(-3'sd3)}}&((3'd5)==(-4'sd7))));
  localparam [5:0] p2 = (-(&(~(({2{(5'sd12)}}^~(^(2'd2)))===((-3'sd3)<<(3'sd1))))));
  localparam signed [3:0] p3 = ((((5'd22)<<<(5'd13))==((3'sd3)===(-4'sd1)))|(((2'sd1)|(5'd8))-((5'd24)<=(2'd2))));
  localparam signed [4:0] p4 = (4'd2 * ((2'd2)?(2'd2):(5'd10)));
  localparam signed [5:0] p5 = {2{(~|(((4'sd5)?(4'd10):(5'sd15))?((-2'sd0)?(5'sd12):(-2'sd0)):(&(5'd13))))}};
  localparam [3:0] p6 = ({4{(+(-3'sd2))}}+(|(((3'd4)&&(-4'sd2))?{(3'd5)}:((3'sd0)?(2'sd0):(5'sd2)))));
  localparam [4:0] p7 = (-4'sd0);
  localparam [5:0] p8 = {1{{1{((4'd12)+({4{(-5'sd9)}}&{4{(5'sd10)}}))}}}};
  localparam signed [3:0] p9 = {((2'd1)>(2'd1))};
  localparam signed [4:0] p10 = {(((4'd10)<(4'd8))&((-2'sd0)+(5'd30)))};
  localparam signed [5:0] p11 = {{{(5'sd13),(-3'sd0),(4'd15)},{(2'sd1),(3'd6)}},{(-2'sd0),(4'd13),(2'sd1)}};
  localparam [3:0] p12 = (3'd5);
  localparam [4:0] p13 = ((3'd2)^~(2'sd1));
  localparam [5:0] p14 = (~({(|(5'sd0)),{(2'd1),(3'sd2)}}?((4'd2 * (4'd15))>>((-2'sd0)?(3'd6):(5'd24))):(~|((2'd3)&&(5'd5)))));
  localparam signed [3:0] p15 = {2{(~|({1{((5'd22)<<(3'd1))}}<=((-3'sd0)>>>(4'sd5))))}};
  localparam signed [4:0] p16 = (2'd3);
  localparam signed [5:0] p17 = ({((~&{2{(-5'sd10)}})!={(3'sd1),(5'sd4),(4'd0)})}>>{{{(4'd4)}},{(5'sd4)}});

  assign y0 = {1{{1{(2'd2)}}}};
  assign y1 = (^((^(p17?p4:p8))?((-p16)+(p5>>p4)):(-(p9?p1:p17))));
  assign y2 = (2'd0);
  assign y3 = (-(((p4?a4:p0)&&(b0?p3:p13))?((!(p6?a5:p10))&&(p2<p1)):((p12?p13:p16)>=(p6/p16))));
  assign y4 = (|(+$unsigned((!(~|a5)))));
  assign y5 = $signed($unsigned($unsigned(((^(~^(&a4)))===(a4?b4:b5)))));
  assign y6 = $signed((($unsigned(b2)<<(a5===a2))>={3{a0}}));
  assign y7 = (-((2'd3)<=(p17?p4:p12)));
  assign y8 = ((-(4'sd4))|{p17,p3,p0});
  assign y9 = {{b1,a0,p6},{p5,p2,a4}};
  assign y10 = {(!p8)};
  assign y11 = (((2'd3)==$signed((a2>>>b5))));
  assign y12 = ((!(a2/a2))>((b1?a5:a5)>>>(a5>>b5)));
  assign y13 = (&(|{4{{2{p9}}}}));
  assign y14 = (-5'sd4);
  assign y15 = (-4'sd6);
  assign y16 = {(+p2)};
  assign y17 = (((a3!==a3)<<(p4>=p9))-{2{(p9?p5:p11)}});
endmodule
