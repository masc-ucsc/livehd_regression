module expression_00922(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((-2'sd1)>(4'd12))==((4'd13)<=(3'd5)));
  localparam [4:0] p1 = {2{{3{((5'd28)?(4'sd6):(2'd0))}}}};
  localparam [5:0] p2 = ((((5'd11)>(3'sd1))<=((4'd9)===(-4'sd1)))&(((2'd1)*(2'd0))*((4'sd5)==(3'sd0))));
  localparam signed [3:0] p3 = (4'd2 * (^(5'd4)));
  localparam signed [4:0] p4 = {1{{3{(((4'd12)===(4'sd5))<<<{1{(4'sd7)}})}}}};
  localparam signed [5:0] p5 = ((~|((3'd3)|(5'd14)))?(((-4'sd6)|(2'sd1))<<((5'd23)^~(3'd1))):((+(2'sd0))==(-(4'd13))));
  localparam [3:0] p6 = (^(2'sd0));
  localparam [4:0] p7 = {4{{2{{4{(4'd11)}}}}}};
  localparam [5:0] p8 = (+(((5'd6)>(5'd7))>>>(5'd11)));
  localparam signed [3:0] p9 = (5'd7);
  localparam signed [4:0] p10 = {{{((4'd10)?(5'd19):(-5'sd4)),{(-3'sd1)},(-2'sd0)},(-4'sd2)}};
  localparam signed [5:0] p11 = {{(-3'sd3),(4'd14),(2'sd0)}};
  localparam [3:0] p12 = ((4'sd1)&(2'd0));
  localparam [4:0] p13 = (&{((5'sd0)||(2'sd0)),{(5'd30),(2'sd0)},((2'sd1)==(3'sd0))});
  localparam [5:0] p14 = ((((-3'sd2)>(-5'sd4))||(|(5'd12)))>>>((~(-3'sd3))!==((4'sd5)<(4'd14))));
  localparam signed [3:0] p15 = ((~{((5'd20)==(-5'sd14)),((2'd0)?(-5'sd7):(2'sd0)),{(3'd0),(3'd5)}})^~{((2'sd1)>>>(4'd1)),((2'd1)?(3'd5):(2'd0))});
  localparam signed [4:0] p16 = {4{(4'd7)}};
  localparam signed [5:0] p17 = (((4'd0)?(2'd2):(2'd0))?((4'd4)?(-5'sd11):(4'd15)):(|((5'd22)?(4'd7):(-2'sd0))));

  assign y0 = (~&(-(4'd15)));
  assign y1 = {(a2>>>a2),(a0+b1),{b3,b2}};
  assign y2 = {2{$signed((|{4{p13}}))}};
  assign y3 = (&($signed($unsigned((!(~((a0!==b2)|(~^a5))))))||((+$signed((|a5)))!=(&(p12&b3)))));
  assign y4 = (4'd14);
  assign y5 = $unsigned((~|({4{p10}}?(p1<<<b2):(+p5))));
  assign y6 = {(p4&&p6),(p13?p1:p4)};
  assign y7 = (~(2'sd1));
  assign y8 = {4{(~|(~(~a3)))}};
  assign y9 = $unsigned((!({4{(|a2)}}&{1{(!{2{{1{a2}}}})}})));
  assign y10 = (4'sd2);
  assign y11 = (a5?p5:p6);
  assign y12 = {2{p8}};
  assign y13 = ((b0?p15:b2)?(4'sd0):(-2'sd1));
  assign y14 = (-4'sd0);
  assign y15 = {4{((a3>>>a0)<<{1{a3}})}};
  assign y16 = $unsigned($unsigned((&$signed((|(-(~^a3)))))));
  assign y17 = $signed(((a4<a3)!==(b0<<<b2)));
endmodule
