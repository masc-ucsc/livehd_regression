module expression_00769(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd5)?(2'd0):(3'd6));
  localparam [4:0] p1 = (-((2'd2)?(-3'sd3):(4'sd5)));
  localparam [5:0] p2 = (&(((4'd10)?(3'sd3):(-5'sd3))?(^(5'sd8)):(~(4'd5))));
  localparam signed [3:0] p3 = ((((5'd23)?(2'd1):(2'sd1))>={(2'd2)})+{3{{3{(2'sd1)}}}});
  localparam signed [4:0] p4 = (-4'sd1);
  localparam signed [5:0] p5 = (+{4{((3'd4)?(5'd30):(-3'sd0))}});
  localparam [3:0] p6 = ({2{((-5'sd2)<<<(3'sd3))}}?({(-3'sd1),(4'sd5)}!=((2'd1)?(5'd0):(3'sd1))):((-5'sd15)?(-4'sd7):(-4'sd1)));
  localparam [4:0] p7 = {{(-2'sd0),((5'sd8)?(3'sd0):(-2'sd0)),((4'd6)>>>(4'd7))},(((2'd0)?(5'd27):(-5'sd6))?(4'd1):{(4'd6),(2'sd1)})};
  localparam [5:0] p8 = (-3'sd2);
  localparam signed [3:0] p9 = ((3'd5)<=(3'sd1));
  localparam signed [4:0] p10 = (4'd12);
  localparam signed [5:0] p11 = {({(5'd4),(3'd7),(4'sd3)}?((3'd4)?(-2'sd0):(5'd13)):{(5'd15),(4'sd1)})};
  localparam [3:0] p12 = (&(&(|(~^(+(|{(((3'd0)>>(5'sd7))+(!(~&(4'sd7))))}))))));
  localparam [4:0] p13 = (3'sd2);
  localparam [5:0] p14 = ((((5'd25)^(2'd3))!==((2'd1)===(4'd6)))<=((4'd2 * (4'd9))<<<(!(3'd5))));
  localparam signed [3:0] p15 = (^(4'd4));
  localparam signed [4:0] p16 = (-5'sd15);
  localparam signed [5:0] p17 = (~^{3{(!((2'sd1)<<<(2'd3)))}});

  assign y0 = (2'sd1);
  assign y1 = {4{{2{p3}}}};
  assign y2 = (&{2{{1{((|a1)?(3'd4):{4{a2}})}}}});
  assign y3 = (((5'd2 * p8)?((p17?p3:p13)):(b5&b5))<(({3{b1}}?(-a2):(a1^a4))^~(!({4{p0}}|(p15==p3)))));
  assign y4 = $unsigned((((b0!=a3)||$unsigned($signed(a4)))<<<(-4'sd1)));
  assign y5 = $signed($unsigned($unsigned(($signed((&(~(&(a3)))))))));
  assign y6 = {2{{3{p4}}}};
  assign y7 = (p16?b1:p1);
  assign y8 = (2'd1);
  assign y9 = ((3'd6));
  assign y10 = {1{{4{({3{b4}}-{3{p4}})}}}};
  assign y11 = (({a3,b5,b3}>={(a4^~b1)})<={(b3>=a3),(a0-b3),{b1}});
  assign y12 = (($unsigned($unsigned(((!p7)^(p12!=p7)))))<=(((-(b5>b3)))===((b2>>a2))));
  assign y13 = (^(($unsigned((a0||b1))==={3{a0}})||{4{{4{a1}}}}));
  assign y14 = (({1{(~{3{p12}})}}|{2{(+p14)}})^~(((a0>b0)!=(p13>>p16))>=(!(+(a0+p13)))));
  assign y15 = (~^(-(|(2'd2))));
  assign y16 = ((~&({p5}?(2'sd1):(a0?b0:a1)))<(|{(~&b5),(~^b4),(a3===b0)}));
  assign y17 = (5'd15);
endmodule
