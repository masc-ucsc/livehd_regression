module expression_00297(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd3);
  localparam [4:0] p1 = {{1{(((4'sd6)^(2'd2))>(3'd3))}}};
  localparam [5:0] p2 = (+((((3'd0)?(-3'sd0):(3'd3))>>>((4'd13)!=(-3'sd3)))>>>{4{(4'd1)}}));
  localparam signed [3:0] p3 = ((5'sd8)&(5'd24));
  localparam signed [4:0] p4 = (5'sd7);
  localparam signed [5:0] p5 = (4'sd7);
  localparam [3:0] p6 = (((4'd6)?(3'd7):(-3'sd2))?((3'sd2)?(5'd24):(-4'sd2)):(3'd2));
  localparam [4:0] p7 = (|{(~(-(2'd1))),{(5'd10),(4'd15),(-4'sd6)},{3{(5'd26)}}});
  localparam [5:0] p8 = (~|{1{(-(&(+(^(4'd12)))))}});
  localparam signed [3:0] p9 = (({(-3'sd0),(4'sd3),(2'sd0)}^~(~&((2'd1)!=(3'sd2))))-(((-4'sd3)?(4'd13):(2'd0))?((-5'sd4)==(2'd3)):(+(4'd7))));
  localparam signed [4:0] p10 = ((((2'd2)<<(3'd3))<{2{(5'sd14)}})>>(|(((4'd6)<<<(-3'sd0))>{3{(-4'sd3)}})));
  localparam signed [5:0] p11 = ((2'd0)||{(5'd2 * (2'd2)),(&(3'sd3))});
  localparam [3:0] p12 = (~^(({2{(4'd3)}}<<<((5'sd4)>>(4'sd0)))-{({(-5'sd12),(3'd1)}^~{(4'd0)})}));
  localparam [4:0] p13 = ((&(5'sd15))>>(~|(2'sd0)));
  localparam [5:0] p14 = ((((3'sd1)?(4'd10):(3'd5))-((4'd2)>(5'sd14)))===(((3'sd3)>(2'sd1))||((-5'sd11)<<<(3'd6))));
  localparam signed [3:0] p15 = (!((-5'sd4)<{((5'd26)^(4'd7)),(~^(-4'sd4)),(~^(2'd3))}));
  localparam signed [4:0] p16 = {2{((+(5'd12))&(-(-2'sd1)))}};
  localparam signed [5:0] p17 = (5'd0);

  assign y0 = ((4'd0)?$signed((p6?p14:p4)):$unsigned((p9?p4:p13)));
  assign y1 = (b2>>b2);
  assign y2 = {3{(~&((p3&&a2)<=(2'sd0)))}};
  assign y3 = $signed({{(b4)},(&(b4?a4:b0))});
  assign y4 = $unsigned((((&{a0,b3,a4}))===(+(|(~&a5)))));
  assign y5 = (5'd2 * (~(!p6)));
  assign y6 = ((a2>>>b2)/p8);
  assign y7 = {{{{(!{{{a1,p14,p0}}})}},(^(~|(~&(+(~&{b0,p5})))))}};
  assign y8 = ((p14?p13:b5)?(p10?p14:a2):{2{p15}});
  assign y9 = {3{$unsigned((p9||p15))}};
  assign y10 = (~&($unsigned((a2||b5))===(a4===b1)));
  assign y11 = ((p13<p10)<<<{a4});
  assign y12 = (^{(~|{p5,b4,b0}),{(p7!=b1),(~^p13)}});
  assign y13 = (&(&{4{(~^$unsigned(a1))}}));
  assign y14 = ((p11<<p12)|(-2'sd1));
  assign y15 = ({p8,p11}!=(-(~|p5)));
  assign y16 = {(~|(4'sd3))};
  assign y17 = (p5+p11);
endmodule
