module expression_00677(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-2'sd1);
  localparam [4:0] p1 = (-(-(((~|(-2'sd1))>>>(5'd2 * (2'd2)))^~(~^((4'sd3)?(3'd5):(4'd6))))));
  localparam [5:0] p2 = ((({4{(2'sd1)}}^~((5'sd11)<<<(3'd4)))>(5'd2 * ((2'd3)>(2'd1))))-(({3{(-2'sd0)}}-{3{(-3'sd2)}})+(((-2'sd1)<<<(3'sd1))^~((4'd11)+(3'd6)))));
  localparam signed [3:0] p3 = (+{3{(5'd25)}});
  localparam signed [4:0] p4 = ((|(((2'd3)<(4'd7))<<<(!(2'sd1))))<=(~&(((3'd4)<=(-3'sd3))^~(2'd2))));
  localparam signed [5:0] p5 = (+({{(-4'sd4),(3'sd0)}}<{((5'd31)?(2'sd0):(-4'sd1))}));
  localparam [3:0] p6 = {1{{((5'd18)===(-2'sd1)),((2'sd0)||(3'd2))}}};
  localparam [4:0] p7 = (5'sd0);
  localparam [5:0] p8 = (+({2{(4'd4)}}&&((4'sd0)-(-3'sd3))));
  localparam signed [3:0] p9 = ({1{{3{(4'd14)}}}}<({3{(3'd2)}}==((5'd9)>=(4'd3))));
  localparam signed [4:0] p10 = ((2'sd1)?((3'sd1)&&(5'd28)):((3'd1)?(4'd10):(4'sd1)));
  localparam signed [5:0] p11 = ((((-5'sd4)>>(4'sd2))?((2'sd1)!==(-2'sd0)):(~|(2'd0)))<=((&(3'd0))?((2'd2)?(5'sd7):(-2'sd0)):((2'sd1)-(4'sd0))));
  localparam [3:0] p12 = (4'd11);
  localparam [4:0] p13 = (2'd3);
  localparam [5:0] p14 = {2{(5'sd3)}};
  localparam signed [3:0] p15 = {3{((2'sd1)<=(3'sd0))}};
  localparam signed [4:0] p16 = ((+((4'd3)!=(2'sd1)))&&(^((5'sd10)&(4'sd1))));
  localparam signed [5:0] p17 = (~|(~&(((2'd1)?(2'd2):(-5'sd12))?(((2'd0)?(4'sd6):(-3'sd2))<<(+(-2'sd0))):((~^(-3'sd0))*((4'd9)<(-3'sd0))))));

  assign y0 = (~(-3'sd3));
  assign y1 = ((((p17^~p10)<<(p12|p1))^~((3'sd1)>(-4'sd5)))==(((p3*p4)^(3'sd2))&&(4'd7)));
  assign y2 = (((~p14)?(-p10):(a0?p17:p12))^~((&p6)?{a5,p15}:(p13==p0)));
  assign y3 = (~&(((a0?a5:b1)!=={2{a1}})&{2{(2'd3)}}));
  assign y4 = (-5'sd10);
  assign y5 = ((p17?p2:p5)+(!(p6|p10)));
  assign y6 = {2{((+p4)?(|p8):(~^p9))}};
  assign y7 = (4'd9);
  assign y8 = ((2'd2)^((b2==a2)>>>(2'd1)));
  assign y9 = ((~((p12?p0:p11)?(^a2):(p3?p10:p7)))?$unsigned((~((&(!p17))))):((a1?p15:p1)?(p16?p3:b2):$signed(p0)));
  assign y10 = ((b1<<b5)<<$unsigned(p4));
  assign y11 = ((+{$signed((~(!p15))),(|(~^(+a3)))})>(~^(~&(~&((b4>>p13)-(~^{a1,a3}))))));
  assign y12 = ((5'd4)<=(~(2'd3)));
  assign y13 = ((((p14?a1:p15)^~(p0?b2:p12))-(a5?b0:a3))>=((+(|(a1&a3)))>>>(|(a4||b1))));
  assign y14 = ((p2!=b0)/a0);
  assign y15 = (-5'sd5);
  assign y16 = (4'd2 * (b1^a0));
  assign y17 = (((b1*b4)&(!(b4)))+((2'd0)<<$unsigned((p3))));
endmodule
