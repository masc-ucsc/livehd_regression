module expression_00620(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~|(((3'sd1)<=(4'd4))>>((3'd5)>=(2'sd1))));
  localparam [4:0] p1 = ({3{(-5'sd1)}}||{1{{{3{(-2'sd1)}}}}});
  localparam [5:0] p2 = (-(~&{1{(~(-2'sd1))}}));
  localparam signed [3:0] p3 = ((6'd2 * ((3'd0)?(5'd23):(3'd0)))?((5'd26)?(4'sd5):(2'd1)):((-(3'd1))&&(~&(2'sd1))));
  localparam signed [4:0] p4 = (-5'sd14);
  localparam signed [5:0] p5 = ((((-4'sd1)<=(-4'sd7))+((-3'sd1)!=(-4'sd5)))?(-(((-3'sd1)?(3'd4):(-3'sd1))-((3'd0)===(3'd5)))):(|((-2'sd0)?(2'd2):(4'sd2))));
  localparam [3:0] p6 = {2{{2{{3{(-2'sd1)}}}}}};
  localparam [4:0] p7 = ({4{(5'd8)}}<<{2{(-5'sd3)}});
  localparam [5:0] p8 = {(+{(5'd12),(-2'sd1)}),{(3'sd2),(2'd2),(-2'sd0)}};
  localparam signed [3:0] p9 = {{(~^{{4{(2'd1)}}})},(~^{(^(!(-4'sd7)))}),(~&(~^(!{3{(-4'sd1)}})))};
  localparam signed [4:0] p10 = (^{(3'd3),(-2'sd0)});
  localparam signed [5:0] p11 = {(~|(((5'd29)===(5'd29))-((-4'sd6)==(3'sd3)))),((-4'sd0)>((-3'sd0)-(4'sd2))),{2{{(4'sd7),(4'd1)}}}};
  localparam [3:0] p12 = ((3'd1)=={3{(-3'sd1)}});
  localparam [4:0] p13 = ({2{{4{(-3'sd2)}}}}^~((!(5'd0))==(-(3'd1))));
  localparam [5:0] p14 = {{((-4'sd0)?(-2'sd1):(4'sd3)),((-4'sd5)?(-3'sd0):(5'd26)),((3'sd3)^~(2'sd1))}};
  localparam signed [3:0] p15 = ((((2'd1)>(3'sd1))<((3'sd3)?(5'sd11):(3'd6)))===(((5'd2)>>(2'sd0))?{(4'd13),(-5'sd10),(2'd2)}:{(3'd4),(-2'sd0)}));
  localparam signed [4:0] p16 = {4{{3{(4'sd7)}}}};
  localparam signed [5:0] p17 = ((5'd21)-(2'sd1));

  assign y0 = (&((((&{4{p14}})^{3{p10}})==(^(-$unsigned(((b4===b5)>>>$signed(p14))))))));
  assign y1 = (p9<<<a2);
  assign y2 = ((~|(~&(5'sd9)))-(($unsigned(b3)+(p17<<<p2))>(!(~(+a5)))));
  assign y3 = ({(-(+b1)),(+(-a0))}>={(~(~|b5)),((~|p0))});
  assign y4 = (4'd2 * (!(p12|b1)));
  assign y5 = {3{{4{p7}}}};
  assign y6 = {((+(&$unsigned(p13)))<=((b5<p6)-(b3!==b0))),{{2{(p8|a1)}},{a2,p11,p0}}};
  assign y7 = (-(3'sd0));
  assign y8 = (^(((~^(a4<<<p11))<=(|(!b0)))^~(-((&(~&b2))&(b2?a3:b2)))));
  assign y9 = (((p11?p5:b2)>(a4?p0:p14))<<<($unsigned($signed($unsigned($signed(p5))))));
  assign y10 = ((!(a5===b1))%p8);
  assign y11 = (5'd30);
  assign y12 = ((-(-4'sd5))>(-5'sd0));
  assign y13 = ((-(&(b2!=b5)))?(((a2^~b4)||(~^p0))):$unsigned($signed((p9?p17:p12))));
  assign y14 = (3'sd1);
  assign y15 = (4'd11);
  assign y16 = {{({p17}=={4{p1}}),{{4{b2}}}},$signed(((b1===a1)>(p15>>p4)))};
  assign y17 = ({2{{$unsigned(a3),(b5>=b4)}}}<{2{(~^{1{{a0}}})}});
endmodule
