module expression_00395(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~(((-2'sd1)|(4'sd1))<=((-5'sd7)/(-5'sd15))))||(3'd1));
  localparam [4:0] p1 = (~^((3'd4)^~(-3'sd0)));
  localparam [5:0] p2 = ((!{3{(5'd29)}})=={3{{(2'd3)}}});
  localparam signed [3:0] p3 = (((3'd1)&{2{(2'd3)}})==={3{(-2'sd0)}});
  localparam signed [4:0] p4 = ((((4'd12)<<(5'd4))<={(-2'sd0),(-4'sd7),(4'sd7)})>>>(-2'sd1));
  localparam signed [5:0] p5 = ((~^(-(|((3'sd0)>=(3'd6)))))<<({(2'sd0),(2'sd1),(-2'sd0)}>>(^(!(3'd6)))));
  localparam [3:0] p6 = ((((2'd3)===(-4'sd1))<((-5'sd11)||(3'd0)))||((5'sd8)<<((-3'sd2)>=(4'd6))));
  localparam [4:0] p7 = (!(((3'd1)?(2'd3):(5'd12))&(|(~|(-(2'sd1))))));
  localparam [5:0] p8 = ({1{(4'd11)}}?{2{(3'sd3)}}:((3'd7)?(-3'sd3):(4'sd0)));
  localparam signed [3:0] p9 = ((-(&(((-3'sd0)^~(2'd0))<<<((2'd2)<(5'sd1)))))<=((((4'd12)>=(4'd6))/(3'd3))&(((2'd2)<(4'd11))==((-3'sd0)|(4'sd2)))));
  localparam signed [4:0] p10 = (2'sd0);
  localparam signed [5:0] p11 = {((5'd8)?(-4'sd5):(-4'sd4))};
  localparam [3:0] p12 = (~{(-5'sd12)});
  localparam [4:0] p13 = (((-4'sd4)!==(2'd2))/(4'sd1));
  localparam [5:0] p14 = (~(&(+((-2'sd0)-(2'sd1)))));
  localparam signed [3:0] p15 = (((-3'sd3)^~(+(2'd0)))^~(((-5'sd10)?(4'd13):(5'd13))>((5'd17)!==(3'd1))));
  localparam signed [4:0] p16 = {{((5'd23)&&(3'd6)),(+(3'sd3)),{(4'sd4)}}};
  localparam signed [5:0] p17 = ((+(3'sd2))?((2'd3)===(2'd3)):(~(-4'sd3)));

  assign y0 = (~$unsigned({((a2>a5)!=(b4>a1)),(((a3<a2)-$signed(b5))),{(b1||a2),{b5,b3,b3},{b5,b3}}}));
  assign y1 = (p0==b4);
  assign y2 = {{2{(6'd2 * p13)}},((p4&p13)&{2{p8}}),{4{p15}}};
  assign y3 = $signed($unsigned(((&$signed({2{(p7?p15:p11)}}))?((^($signed(p17)&{1{p7}}))):(+(4'd10)))));
  assign y4 = (({4{b1}}?(b5?b1:a5):{1{(p5>>>a3)}})<<<{2{((-3'sd0)&(5'd21))}});
  assign y5 = ((-((+$unsigned(p8))?(a2>b0):$unsigned((a1>b2))))<<$unsigned((^(5'sd1))));
  assign y6 = (~|(^(((b5)>>(p14?a3:p4))&($unsigned(a1)&&(p9^~p15)))));
  assign y7 = $unsigned(((~&(((p5<=b5)>=(b3>>b3))))>>(|(&((-a5)>={b0,a5,a1})))));
  assign y8 = (^(~^{3{(((|{2{a0}})))}}));
  assign y9 = $signed((5'd29));
  assign y10 = {(-2'sd1),(a4&a1),(a5&a0)};
  assign y11 = $unsigned((p3?b4:p7));
  assign y12 = {4{{2{p12}}}};
  assign y13 = ((-5'sd4)|(((a3*b0)===(a4?b0:b4))+(!(b4-p16))));
  assign y14 = {p8,p11};
  assign y15 = (((b4!==b1)?(b4<=a0):(b1==a1))?(^((-(b3/b3))||((b4/a0)))):(((a2<<a2))===(a3^a1)));
  assign y16 = $signed(($unsigned($unsigned(b0))===(b0-b5)));
  assign y17 = ((a4!==a5)?{p0,p16}:(b5!=p0));
endmodule
