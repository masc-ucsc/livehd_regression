module expression_00397(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((+(|((-5'sd7)&&(-2'sd0))))&(~|((2'd0)>=(2'sd1))));
  localparam [4:0] p1 = ((5'd12)^~(3'd1));
  localparam [5:0] p2 = ((3'd3)?(4'sd4):(-5'sd11));
  localparam signed [3:0] p3 = (^{(^((4'd6)?(2'sd1):(4'd1))),((3'd2)-(2'd0)),((3'sd1)^~(2'd1))});
  localparam signed [4:0] p4 = {1{((2'd0)?(4'd6):(5'd1))}};
  localparam signed [5:0] p5 = ((((5'd5)&(2'sd0))|((2'sd0)&&(-5'sd10)))<={1{((~|(3'sd3))<<(~&((3'sd3)^~(4'd7))))}});
  localparam [3:0] p6 = {{(-{(-5'sd12),(4'd8),(-4'sd6)}),((5'd28)<=(2'd2))},{2{(~&(-(-5'sd4)))}}};
  localparam [4:0] p7 = (((~^((-4'sd0)!=(-5'sd6)))||((2'd3)<=(5'd10)))<((+(&(2'sd0)))^~((2'd1)>=(2'd3))));
  localparam [5:0] p8 = ((((4'd4)+(3'sd3))>((3'd2)^~(2'sd1)))?{3{(5'sd8)}}:{1{{3{(5'sd8)}}}});
  localparam signed [3:0] p9 = {((5'd24)!==(4'sd0)),((3'd0)<(5'd5)),{(-5'sd8),(2'sd0),(4'sd2)}};
  localparam signed [4:0] p10 = {(3'sd3),((~(5'd3))|(-3'sd0)),((5'd10)>=(5'd26))};
  localparam signed [5:0] p11 = ((4'sd1)|((4'sd3)==(3'd2)));
  localparam [3:0] p12 = ((3'd7)?(-3'sd0):(5'sd10));
  localparam [4:0] p13 = (2'd3);
  localparam [5:0] p14 = (~({(3'd2),(!(4'd1)),(5'd22)}+(-(4'd2 * (~^((3'd0)===(4'd11)))))));
  localparam signed [3:0] p15 = ((4'd4)<<(3'd6));
  localparam signed [4:0] p16 = ({((4'sd6)&&(2'sd1))}?{1{((5'd18)?(3'sd2):(5'd27))}}:{4{(3'd1)}});
  localparam signed [5:0] p17 = (-(((-(-5'sd12))>=((2'd3)?(-4'sd3):(-5'sd8)))?((3'd2)?(2'sd0):(2'd3)):((&(3'd0))||((5'd31)?(-2'sd1):(2'd0)))));

  assign y0 = (a2?p13:p3);
  assign y1 = (~{2{((a5^~p13)==(+a2))}});
  assign y2 = ({2{b4}}<<{4{a0}});
  assign y3 = (^((b1*p2)==(a5%a5)));
  assign y4 = (-5'sd6);
  assign y5 = ($signed(((b4<<a4)==(a4?b2:a4)))<<<({1{(a4?b2:a2)}}==(b4?a4:a5)));
  assign y6 = ({a0,b4,a5}&(b1>b4));
  assign y7 = (2'd1);
  assign y8 = {2{$signed($unsigned(({a5,a1,b1}!==(b2?a2:b5))))}};
  assign y9 = {{1{{3{(-2'sd0)}}}}};
  assign y10 = (~{((-4'sd5)),(~|((4'd11)-(4'sd5)))});
  assign y11 = $unsigned((({3{b3}}===(b1<<b1))<={4{a5}}));
  assign y12 = ((-3'sd0)>>(~|$signed((p16!=p13))));
  assign y13 = ((a5&&a2)^$signed((~|b0)));
  assign y14 = $unsigned({3{(p1-a4)}});
  assign y15 = (~&((~|((b4?a2:a3)===((a2^~a2))))&((p6>=a2)?(p15<<<a4):$unsigned((5'sd6)))));
  assign y16 = {((a2||b1)==(b0>=b4))};
  assign y17 = ((+(($unsigned((^b2))^~(p0<=p1))^~$unsigned((~^(((~p17))/p1))))));
endmodule
