module expression_00774(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (5'd2 * ((2'd1)&&(3'd2)));
  localparam [4:0] p1 = (~^(~^(3'd3)));
  localparam [5:0] p2 = (~(-4'sd7));
  localparam signed [3:0] p3 = ((&(~(-5'sd6)))?(-2'sd1):((2'sd0)?(5'd20):(4'd0)));
  localparam signed [4:0] p4 = (((&(4'sd5))?((2'd3)?(2'd0):(2'd0)):((2'd2)>>(3'd0)))?(-((~^(2'sd0))!=={(-3'sd2),(3'd6),(3'd5)})):(|((-3'sd1)?(-5'sd9):(5'd16))));
  localparam signed [5:0] p5 = (!(+((((-4'sd5)?(3'd0):(5'd21))<<<(~&(4'sd2)))?((2'd3)?(-3'sd2):(4'd0)):((3'sd0)?(4'd5):(5'sd9)))));
  localparam [3:0] p6 = {3{(3'd5)}};
  localparam [4:0] p7 = (&(((5'd19)?(-3'sd1):(3'd0))?(5'sd10):(!((5'sd9)?(-3'sd2):(3'd6)))));
  localparam [5:0] p8 = (((((5'd5)/(3'sd3))^(&(5'd13)))^~(~(-(~(2'd0)))))>((^(&((3'sd0)%(-2'sd0))))+(((3'd5)!==(2'sd1))<<(+(-3'sd3)))));
  localparam signed [3:0] p9 = (3'sd3);
  localparam signed [4:0] p10 = (~&(((2'd0)>>>(4'd12))/(2'd2)));
  localparam signed [5:0] p11 = (((((5'd30)^(4'd15))>>>((-2'sd0)?(-2'sd1):(2'd2)))&&(^(~|((3'sd0)?(4'd2):(-3'sd0)))))^(((3'd5)>(4'sd0))?((5'd13)?(4'sd4):(-3'sd0)):((5'd17)?(3'd1):(4'd15))));
  localparam [3:0] p12 = {2{(-4'sd0)}};
  localparam [4:0] p13 = ((4'd2 * ((5'd12)^(5'd19)))<(4'd2 * ((3'd4)!=(4'd5))));
  localparam [5:0] p14 = ((!(~(4'd8)))<=(|((2'sd0)&&(4'sd0))));
  localparam signed [3:0] p15 = {4{{{(-4'sd2)}}}};
  localparam signed [4:0] p16 = (5'd2 * {(4'd15),(3'd7)});
  localparam signed [5:0] p17 = {2{(((3'sd0)^(4'd12))^~((2'd1)^(5'd23)))}};

  assign y0 = (!$signed((~^(~|(|(p1?p0:p5))))));
  assign y1 = {(4'd2 * p1),(&(b0?p3:p14))};
  assign y2 = ($unsigned((~^$signed({p12,p17,p11})))?($unsigned((p8?p2:p0))>>>{(a0?p10:p8)}):{({p8,p5}||(b3?p10:p13))});
  assign y3 = (((p15?b1:a0)>(p6?a1:p12))?({b5}&&(b4+a1)):({4{a5}}>>(4'd2 * a0)));
  assign y4 = ((((-(!(|$unsigned((-b5)))))|(~$unsigned((~&((a3!=b1))))))));
  assign y5 = {((2'd1)-(p5>>>p4)),(2'd0),((6'd2 * p2)!=(p13||p11))};
  assign y6 = (+(((~&(|(+a1)))&((~|a4)<<(~a4)))===((&(~^(a5>>>a0)))<<(6'd2 * (a0!==b0)))));
  assign y7 = ((5'd2 * {4{a1}})!=={4{{3{a0}}}});
  assign y8 = ((a2?p15:b4)<(~&(b5<p13)));
  assign y9 = ((4'd4)?(5'sd6):{{a4,a4},{a2,a1,a3}});
  assign y10 = (($signed((p17))<=(a5>>>p12))<((~&(p3>>>p9))^~(p10<=a4)));
  assign y11 = {2{(~&{1{({1{{4{b2}}}})}})}};
  assign y12 = (b1&&a4);
  assign y13 = (2'd0);
  assign y14 = ((~&p10)^{p12,p10,p7});
  assign y15 = {2{(5'd31)}};
  assign y16 = (-(~|$unsigned($signed({3{((p7+p10)!=(+(b5!==b1)))}}))));
  assign y17 = $signed($signed((p8&&p6)));
endmodule
