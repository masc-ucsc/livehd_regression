module expression_00927(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-(((3'sd2)-(-2'sd0))>=(~&(4'd9))));
  localparam [4:0] p1 = ((-3'sd2)!=={(3'd0),(2'd2)});
  localparam [5:0] p2 = (~&((&(!(4'd2)))>>>((-4'sd6)<<<(-3'sd2))));
  localparam signed [3:0] p3 = {{(~^(!(!((5'sd7)===(-5'sd14))))),(-4'sd5),{((-5'sd1)|(-3'sd2)),(~|(2'sd1))}}};
  localparam signed [4:0] p4 = (!({(5'sd10),(4'd1),(4'sd3)}||((5'd14)<(-2'sd1))));
  localparam signed [5:0] p5 = (3'd5);
  localparam [3:0] p6 = ((-2'sd1)^(((3'd3)%(5'sd10))==((2'sd0)+(3'd1))));
  localparam [4:0] p7 = (~|((-2'sd1)||(2'sd1)));
  localparam [5:0] p8 = (((3'sd0)?(2'd2):(5'd27))?(2'd3):(-5'sd9));
  localparam signed [3:0] p9 = (4'd5);
  localparam signed [4:0] p10 = (3'sd1);
  localparam signed [5:0] p11 = ((((2'sd1)-(5'd21))<<<((4'd10)!=(4'sd4)))!==({(-4'sd2),(4'sd0),(5'sd13)}&((4'sd3)&(-2'sd0))));
  localparam [3:0] p12 = {2{({1{(+{2{(2'sd1)}})}}-{4{(2'sd1)}})}};
  localparam [4:0] p13 = (5'sd11);
  localparam [5:0] p14 = (|(3'd7));
  localparam signed [3:0] p15 = ((((4'd11)?(3'd3):(2'd2))?((5'd22)?(2'd1):(-4'sd1)):{4{(5'sd0)}})?(((5'sd0)?(5'sd11):(-3'sd0))?((5'sd7)?(5'd18):(2'd2)):(-(4'd0))):{2{(^(-3'sd3))}});
  localparam signed [4:0] p16 = ({((5'd5)+(3'd4))}&((-2'sd1)^~(5'sd11)));
  localparam signed [5:0] p17 = {((+(5'sd8))<<<{(2'sd0),(3'd5)}),(-{{(5'd15),(-2'sd0),(-3'sd2)}}),{(2'd0),(5'd0),(4'd9)}};

  assign y0 = ((~^$unsigned((~|((&a4)&&{p9,p1,p1}))))>>>{(b1-b0),(-p16),(p5^~p12)});
  assign y1 = {a2};
  assign y2 = (((4'd12)?(b1-p6):(p3&&a1))<<(|((a2?p12:p8)?(a3?p16:a5):(p14?p17:a3))));
  assign y3 = {3{{1{p15}}}};
  assign y4 = (-((3'sd0)===((a1+b0)|{4{b3}})));
  assign y5 = ({1{($unsigned($unsigned({3{$signed(a1)}}))||({4{a1}}<{1{{2{b0}}}}))}});
  assign y6 = (~(-((~&{(~a1),(p8>>>b3)}))));
  assign y7 = $signed((({(({b3,b4}<<(a0))===((|a3)<={b3,b5})),(~&(-5'sd15))})));
  assign y8 = (5'd0);
  assign y9 = (((p5>p8)?(&(^p9)):{{3{p9}}})&{2{(3'd2)}});
  assign y10 = ((3'd0)>>>(p11?a2:a3));
  assign y11 = $signed((($unsigned($signed($unsigned(($unsigned(($signed($signed($signed($unsigned($signed(($signed($signed($signed($signed(p4)))))))))))))))))));
  assign y12 = (~(-((~&(4'd3))?(|(~&b1)):(b0?b4:a3))));
  assign y13 = {(-(b0<<<a5)),{b0,a1}};
  assign y14 = {{(b1>a2)},(4'd2 * (b0-p12)),{a1,b5,a3}};
  assign y15 = ({{2{p10}},(a0<<a5),(b0!=a2)}&(2'd2));
  assign y16 = $unsigned((-(&(+{(({a2,p8}&{a1,a2})^~$signed($signed((p6+p16))))}))));
  assign y17 = (&(^(a4?b0:a5)));
endmodule
