module expression_00715(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'd10)!=(4'd15))|(!((4'd9)>>(3'd0))));
  localparam [4:0] p1 = (((5'd0)?(-2'sd1):(-2'sd1))>={2{(+(2'd0))}});
  localparam [5:0] p2 = {1{{1{(2'd3)}}}};
  localparam signed [3:0] p3 = ((|(&(!(5'sd8))))?((-(4'd6))===(~(4'd7))):((-5'sd7)?(-2'sd0):(3'd0)));
  localparam signed [4:0] p4 = ((!((3'sd0)?(3'sd2):(3'sd2)))<=((-2'sd1)?(-2'sd0):(-2'sd1)));
  localparam signed [5:0] p5 = (+(^((((-5'sd0)!=(3'd7))!=={3{(-5'sd4)}})<<<{2{{4{(5'd2)}}}})));
  localparam [3:0] p6 = (2'sd1);
  localparam [4:0] p7 = (~|(((4'sd3)?(5'sd13):(2'sd1))?(-4'sd5):((2'd2)?(-3'sd0):(3'sd2))));
  localparam [5:0] p8 = ((-((2'd0)?(5'sd10):(4'd11)))?((4'd15)?(4'd13):(5'sd1)):(2'd2));
  localparam signed [3:0] p9 = {1{{4{(-(2'd1))}}}};
  localparam signed [4:0] p10 = (&{{((2'sd0)+(2'd1))},((~^(2'sd1))||((2'd0)==(3'sd1))),(~^{(5'd13),(5'sd6),(3'd0)})});
  localparam signed [5:0] p11 = (3'd7);
  localparam [3:0] p12 = ((~&((5'd7)?(3'sd0):(3'sd2)))>>>((-4'sd3)?(5'd31):(2'd0)));
  localparam [4:0] p13 = (((+(-2'sd0))?((2'd0)?(3'sd1):(3'd7)):((3'd0)?(5'd1):(-4'sd2)))-(&(((2'd1)>(2'd3))<<<(-(4'd11)))));
  localparam [5:0] p14 = ((((2'd3)!=(3'd2))?((2'sd1)>=(-3'sd3)):((-3'sd3)?(5'sd14):(5'd7)))?((5'd16)?((2'sd0)-(4'd5)):((-5'sd4)?(5'd13):(2'd0))):(((-3'sd1)<=(2'sd0))<((3'd4)===(2'd3))));
  localparam signed [3:0] p15 = (-{{{(-3'sd0),(-4'sd4),(5'd25)},(~|(+(2'd1)))},(~^{(~|(-3'sd1)),{(-2'sd1),(-2'sd0)},(|(2'd3))})});
  localparam signed [4:0] p16 = ((2'd1)?(5'd19):(2'd3));
  localparam signed [5:0] p17 = (~^(5'd2 * {1{(~(3'd3))}}));

  assign y0 = {1{(~&({2{((p12&&p15)?{1{(p3==a0)}}:(p16<=p14))}}))}};
  assign y1 = (~(((a1===a4)<{1{b5}})?((b5?b0:b2)&{a1,b4}):((b0?b5:a1)?{1{a5}}:{2{p15}})));
  assign y2 = {1{{{((p17&p12)>>(~&(p11&&p13)))},{{2{{1{{2{p1}}}}}}}}}};
  assign y3 = (-(-p4));
  assign y4 = (3'd5);
  assign y5 = {(~(|({4{p0}}==(p10&&p17)))),({4{p2}}>{p5,p6})};
  assign y6 = (a5?b3:p11);
  assign y7 = ((4'd14)^~$signed({(2'd3),{p4,a0,p13}}));
  assign y8 = ((2'd2)?$signed(((p6?p1:p17)?(p4?p4:p1):(p5&&p2))):((p7^a3)/p0));
  assign y9 = $signed($signed((((b5?b5:a4)&(b2?b0:a1))-((a5==a5)?{2{a1}}:(b1>>a3)))));
  assign y10 = (3'sd2);
  assign y11 = (+(~|{(+(^(&{(~|b1)}))),{{p10,p15,p12},(+{b3})},(|{(-a1),(&p5),{p1}})}));
  assign y12 = ((b1>=p12)&{3{p9}});
  assign y13 = $unsigned(((|((b0&&p12)||(~|(b4<<<a0))))==(((5'd30)!=(a1^a4))^~({2{a4}}===(b2)))));
  assign y14 = (({3{b2}}<{(b2!=a0),{b4,p12,b0}})>>>(4'sd0));
  assign y15 = (-((^(-{b5,a5,b3}))!==(b3?a2:b4)));
  assign y16 = ((((b2&&a0)/a5))+($unsigned((-(^(p17<<b5))))));
  assign y17 = (a0^a0);
endmodule
