module expression_00221(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {((3'd5)>>(3'sd3)),{(2'd2),(2'sd1),(-3'sd3)},{(-5'sd7),(3'sd3)}};
  localparam [4:0] p1 = (((5'sd10)>=(2'd0))?((5'd4)?(-3'sd3):(4'sd7)):{4{(4'd1)}});
  localparam [5:0] p2 = (&(((~&(3'd6))>>(|(3'sd2)))<<<{(2'd2),(4'd3),(3'sd3)}));
  localparam signed [3:0] p3 = {{{(4'd10),(3'd3),(5'sd0)},{(-5'sd7),(5'sd12),(5'sd6)},{(2'sd1),(3'sd0)}},{{(4'd2)},{(-3'sd2),(4'd4)},{(3'd0)}}};
  localparam signed [4:0] p4 = {2{((2'sd0)?(4'd9):(3'd2))}};
  localparam signed [5:0] p5 = ((4'd0)<<<(3'd5));
  localparam [3:0] p6 = {3{{2{((2'sd1)?(5'd25):(5'd14))}}}};
  localparam [4:0] p7 = {4{{(~(5'sd13)),((5'd27)<(4'd15))}}};
  localparam [5:0] p8 = ((~&(3'sd0))^~{(+({(5'sd1)}===(2'sd0)))});
  localparam signed [3:0] p9 = (~&(-((2'd2)?(3'd0):(2'sd1))));
  localparam signed [4:0] p10 = {4{{(3'sd2),(2'd2),(5'sd4)}}};
  localparam signed [5:0] p11 = (!{(3'sd0),(2'sd1),(5'd19)});
  localparam [3:0] p12 = (~&(|(^((5'd7)>=(2'd3)))));
  localparam [4:0] p13 = (((-2'sd0)?(5'sd14):(4'd11))?((3'd6)?(3'sd0):(-2'sd1)):(2'd2));
  localparam [5:0] p14 = ({(2'sd1),(3'd6)}?{(5'd28)}:{4{(4'sd0)}});
  localparam signed [3:0] p15 = {2{{2{(2'sd0)}}}};
  localparam signed [4:0] p16 = {4{{2{(3'sd3)}}}};
  localparam signed [5:0] p17 = (&(&(-(^(~|(2'sd1))))));

  assign y0 = (((p1+a2)?{a3,a5,b5}:(p3-b3))?($unsigned((p11>=p1))):((b0^p0)?(p5>>b4):(a1?b0:p7)));
  assign y1 = {(-(2'd3)),(~{(~&b5)})};
  assign y2 = ({({a1,a1}),((b1>=a4))}!==(-4'sd1));
  assign y3 = ((~&((p2?a2:b5)?(-2'sd1):(b4?p13:a0)))?(-2'sd1):(-5'sd12));
  assign y4 = $unsigned((b4?b4:p7));
  assign y5 = (4'd9);
  assign y6 = ({2{$unsigned((+(~^{4{a0}})))}});
  assign y7 = ((((b4)>>(3'sd3))>>((p9>>p9)))||$signed((-5'sd7)));
  assign y8 = {1{b5}};
  assign y9 = ($signed($signed((-4'sd7)))<=$signed((p5?b3:a5)));
  assign y10 = (-4'sd6);
  assign y11 = (((p3==p3)>(p10<p12))^~(-(~&(p13^p14))));
  assign y12 = {4{p7}};
  assign y13 = {1{{{2{({1{b1}}+{a4,b1,a4})}},(((b4!==a2)===(b0>>>a1))+({p4}>{a0,b3}))}}};
  assign y14 = {(p13==p12),$signed(a2)};
  assign y15 = (+(~&(~$signed(((~(~&(p5&p0)))^$signed((~|(5'd2 * p1))))))));
  assign y16 = ((6'd2 * p14)>>{a5,p16});
  assign y17 = {4{(+(-4'sd3))}};
endmodule
