module expression_00717(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd1)?(4'd8):(-2'sd0))<(^((-5'sd3)>(5'd18))));
  localparam [4:0] p1 = ((3'd2)?(-3'sd3):(4'd9));
  localparam [5:0] p2 = ((((-4'sd6)^(2'sd1))/(5'sd14))<(((-3'sd0)+(-3'sd2))>>>((-4'sd7)>>(5'sd2))));
  localparam signed [3:0] p3 = (3'sd3);
  localparam signed [4:0] p4 = ((5'd2 * {2{(2'd0)}})>={(4'd2 * (2'd3))});
  localparam signed [5:0] p5 = (&(4'sd7));
  localparam [3:0] p6 = {1{((&(5'sd5))?{(-3'sd3),(2'd3)}:{(2'd3),(5'sd7)})}};
  localparam [4:0] p7 = {(^(^(+(~|(3'd3))))),(+(&((-4'sd0)-(5'd7)))),(~{((2'd2)<=(5'd11)),(~|(-3'sd1))})};
  localparam [5:0] p8 = {2{(-5'sd3)}};
  localparam signed [3:0] p9 = (~((~^(((5'd4)|(2'sd1))&((-2'sd1)^~(4'd5))))>>(((-2'sd0)&(3'd1))?((4'd12)||(2'd1)):((-5'sd12)>=(-3'sd1)))));
  localparam signed [4:0] p10 = (-2'sd0);
  localparam signed [5:0] p11 = ((+((-4'sd1)?(-2'sd0):(2'd3)))?((|(5'd20))===(&(3'd4))):(((5'sd5)||(-4'sd7))==((5'd0)?(-4'sd2):(2'd2))));
  localparam [3:0] p12 = {3{(((3'sd0)?(2'd2):(5'd28))?{3{(-2'sd1)}}:(&(3'd4)))}};
  localparam [4:0] p13 = {1{(((4'sd4)&(3'd5))==((3'd3)&(-3'sd0)))}};
  localparam [5:0] p14 = {1{(4'd15)}};
  localparam signed [3:0] p15 = {((5'd12)?(2'sd1):(3'd7)),(5'd13),(5'd14)};
  localparam signed [4:0] p16 = (2'd2);
  localparam signed [5:0] p17 = {((4'sd0)<<<((4'sd0)===(2'd3))),(-2'sd1)};

  assign y0 = (^((4'd2)^~(((p7>>>p3)-$signed(p0)))));
  assign y1 = (~&$unsigned((~|(({a1}<<(p16))&(+((~a2)>{b1,b1,p7}))))));
  assign y2 = (((+(&b5))=={3{b0}})^~{1{(~^{2{{2{a2}}}})}});
  assign y3 = {1{$signed(((((p0>p0)&{4{p15}})>($signed(p5)-(4'd2 * b0)))&&(((p11<=b4)<(a1===b4))<$signed((p15<<a2)))))}};
  assign y4 = ((^((a0===b2)-(p8==p12)))?((5'sd1)+(b3?p5:p11)):((-4'sd5)>=(~&p13)));
  assign y5 = (-3'sd3);
  assign y6 = {2{(p12^p15)}};
  assign y7 = (((a0?p6:p15)?(b3?p17:p7):(p9?p5:p13))?((p14?p9:b4)>>>(b4?p15:p4)):{((|a0)>>(|p14))});
  assign y8 = (+((~(p12&&a4))>{p4,a4,p10}));
  assign y9 = ((a2!==a2)^(b1>=a4));
  assign y10 = {3{p7}};
  assign y11 = ((~^(!(((p13?p7:p4)))))?((~&(b0?a0:b2))!==(b3?b4:b5)):((p6?p5:a2)>=(p12<<<b3)));
  assign y12 = (-3'sd1);
  assign y13 = (($unsigned($unsigned($signed($unsigned(((^(b3-p16))&&$signed((p13&&b3)))))))||((~((~|p10)>=$unsigned(p16)))^~(+((^p9)<=(~|p2))))));
  assign y14 = $signed({1{$signed(($signed(((($unsigned(p2)))<<<((4'd14)===(b0!==b4))))>>>{1{(4'd14)}}))}});
  assign y15 = (b3==p14);
  assign y16 = (-(~^((+(!(~|b3)))<(5'sd7))));
  assign y17 = {(b5>=p9)};
endmodule
