module expression_00418(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {({1{(5'd19)}}>{2{(-3'sd2)}}),({2{(2'd0)}}===(4'd7)),{{(5'sd7)},{(-4'sd0),(5'd26)}}};
  localparam [4:0] p1 = (((4'sd3)?(-5'sd4):(5'sd12))>>(|{3{(4'sd2)}}));
  localparam [5:0] p2 = ((-((-4'sd1)^~(-2'sd1)))<<<((2'sd0)?(3'd2):(4'd15)));
  localparam signed [3:0] p3 = {2{(((-2'sd1)?(5'd7):(3'd1))<=(((-2'sd0)&&(5'sd5))<<{3{(-3'sd3)}}))}};
  localparam signed [4:0] p4 = (((-4'sd1)+(-4'sd0))>>{2{(-4'sd4)}});
  localparam signed [5:0] p5 = {{{{(4'sd5),(4'sd0),(-3'sd0)}},{(2'sd1),(5'sd0),(2'sd0)}},{{(2'd3),(5'sd4),(2'sd0)},{(2'd3)},{(2'sd1)}}};
  localparam [3:0] p6 = (~|(~|(|((4'sd2)<=(-3'sd3)))));
  localparam [4:0] p7 = (5'sd9);
  localparam [5:0] p8 = {(4'sd0),((2'd0)<(2'd3)),(5'sd9)};
  localparam signed [3:0] p9 = {1{{1{{{{3{{1{(5'sd0)}}}}},{3{{1{(5'd26)}}}}}}}}};
  localparam signed [4:0] p10 = ({1{({1{(4'd9)}}!==(~(3'sd2)))}}&&{2{{(3'd1),(4'd8)}}});
  localparam signed [5:0] p11 = {{{1{(-3'sd1)}},{4{(-3'sd3)}}},{{3{(-2'sd0)}}},((-2'sd0)?(2'sd1):(2'd0))};
  localparam [3:0] p12 = ((2'sd1)!==(4'd0));
  localparam [4:0] p13 = (-5'sd12);
  localparam [5:0] p14 = (((-2'sd1)<<<(2'd0))!=((3'd3)?(-3'sd2):(2'd3)));
  localparam signed [3:0] p15 = ((-(((5'sd4)!=(5'sd9))+(&((2'sd1)<<<(2'd2)))))>>>({((2'sd0)<(5'd31)),(~(3'd1))}^(((5'd27)&(3'd4))+(~&(5'd27)))));
  localparam signed [4:0] p16 = {({(3'sd2),(3'd3)}<=(5'd2 * (4'd7))),(((5'd18)^(4'd11))==={(5'd20),(5'sd2),(-4'sd5)})};
  localparam signed [5:0] p17 = (~|(~|({(4'sd4),(-3'sd2)}+(5'sd7))));

  assign y0 = {(({{p7,p8,p12},(4'd12)}&((3'd6)?(p6<<p17):(a5>>>p7))))};
  assign y1 = ((a3?b3:a4)<<<(b3?a0:a3));
  assign y2 = (((!((^((a3^~a3)===(a0^a5)))))>$unsigned((~^(4'd2 * $unsigned((p17<<p6)))))));
  assign y3 = ((3'd3)<<<(&((~&{b4,a1,a4})<<(b1-b3))));
  assign y4 = (+(4'sd5));
  assign y5 = (2'd3);
  assign y6 = {3{{(p15?p12:p13),(^p0),(b4!==b5)}}};
  assign y7 = ((p10*p8)^~(p16/p2));
  assign y8 = ({4{b1}}<{1{$unsigned(a4)}});
  assign y9 = ((-5'sd6)?((p16?p7:p15)?(b3==p7):(3'd7)):((p4?p15:b2)?(p17?p9:b3):(4'd14)));
  assign y10 = (-5'sd8);
  assign y11 = (p3>=p14);
  assign y12 = $signed({2{{4{$unsigned(p8)}}}});
  assign y13 = {2{((((-4'sd4)^~(p13==b0)))&&((p8+p0)&&$signed(b3)))}};
  assign y14 = (~|({2{{p9,p6}}}+{$signed({p6,p11,b5})}));
  assign y15 = (~^(&{({2{({1{({p17}>$signed(p0))}})}})}));
  assign y16 = (!((|(~&(~(&((b3%a0)^~(b3<<<p17))))))^(((+b4)<<<(b4<=b3))!=(~(&(~a0))))));
  assign y17 = {((b3?a3:a1)?(p16<<<p15):(b4?a1:b5)),({p11,p2,p11}-(p12<<<p1))};
endmodule
