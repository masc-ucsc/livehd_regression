module expression_00294(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&({(4'sd0),(-3'sd3),(-5'sd4)}?{(5'd26),(5'd31),(-5'sd15)}:(&(-5'sd14))));
  localparam [4:0] p1 = (~(&(2'd1)));
  localparam [5:0] p2 = (((2'd3)?(3'd5):(5'd20))<((-3'sd1)?(-5'sd15):(2'd0)));
  localparam signed [3:0] p3 = ((4'd2 * ((2'd0)-(2'd3)))<<((~|(4'd14))?((4'sd3)?(-2'sd1):(-4'sd2)):((4'sd1)|(-4'sd3))));
  localparam signed [4:0] p4 = (((4'sd2)===(2'd0))&((4'sd0)>(3'd0)));
  localparam signed [5:0] p5 = ((((5'd7)?(5'sd14):(3'd5))+((5'd18)?(4'd1):(-2'sd0)))|(((2'd2)?(2'd1):(-5'sd12))?((5'd15)<<(5'd19)):((5'd0)?(-2'sd1):(2'd1))));
  localparam [3:0] p6 = (-2'sd0);
  localparam [4:0] p7 = {({(-5'sd6),(3'sd1)}+((2'sd1)||(4'd2)))};
  localparam [5:0] p8 = ((((5'd25)>(-2'sd1))>>>((2'd2)^~(-4'sd7)))||(((4'sd1)<=(5'sd1))===(2'sd1)));
  localparam signed [3:0] p9 = {1{(-(~|((4'sd5)-{2{(3'd4)}})))}};
  localparam signed [4:0] p10 = (((3'd2)==(-2'sd0))+((5'd18)<(4'sd0)));
  localparam signed [5:0] p11 = ((6'd2 * (3'd4))*(4'd14));
  localparam [3:0] p12 = (+(((5'd4)||(3'sd2))<<<((-5'sd11)^(4'sd5))));
  localparam [4:0] p13 = ((^((|(4'd3))===((4'd3)===(5'd4))))&(((2'd2)+(-5'sd0))-(6'd2 * (2'd1))));
  localparam [5:0] p14 = ((((-2'sd0)>=(-5'sd14))<=((3'sd3)<<(5'd17)))!=={((-(5'd29))|{(2'd2),(2'd2)})});
  localparam signed [3:0] p15 = (((-2'sd1)<<(2'sd1))==((2'd1)>>(-2'sd1)));
  localparam signed [4:0] p16 = {2{(4'sd4)}};
  localparam signed [5:0] p17 = (+{(4'd3),(4'sd3),(3'd3)});

  assign y0 = (&(~^(~&({3{a3}}>(!b4)))));
  assign y1 = (-(-3'sd1));
  assign y2 = $signed((a3?p6:p17));
  assign y3 = (((^$signed(a0)))===((b0||b5)>$unsigned(a2)));
  assign y4 = (|(-4'sd2));
  assign y5 = ((-3'sd1)>((((5'd1)>>>{2{p14}})!=(2'd0))));
  assign y6 = (|$unsigned((&$signed((((~^(b3+p16))>>>(p13?p2:p6))<<<(+((p9&&p1)>(p17<<<p8))))))));
  assign y7 = (|((3'd3)>>{2{((-p15)>{4{p1}})}}));
  assign y8 = {3{((p1!=p4)<<{4{a4}})}};
  assign y9 = (^(2'd1));
  assign y10 = {{2{(a3-p16)}},((b1^b1)!==(a1?b5:b0)),(-(^(~{3{p16}})))};
  assign y11 = ((~(((~|($unsigned((-3'sd1))))<({(3'd0)}+(p8&&p4))))));
  assign y12 = {3{(-5'sd11)}};
  assign y13 = (~|{4{p0}});
  assign y14 = {(a2?b0:b0)};
  assign y15 = (^(a5?a0:b2));
  assign y16 = $signed({3{{1{{3{p17}}}}}});
  assign y17 = ((4'd15)<<<(4'd9));
endmodule
