module expression_00180(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((2'sd0)?(3'd6):(2'sd1))==(~(4'd6)))===({(4'd7),(3'd0),(3'd4)}||((5'sd0)?(-4'sd3):(3'd0))));
  localparam [4:0] p1 = {4{(-3'sd0)}};
  localparam [5:0] p2 = (6'd2 * ((3'd4)?(3'd4):(5'd17)));
  localparam signed [3:0] p3 = {1{((3'd7)===((4'd0)-(-2'sd1)))}};
  localparam signed [4:0] p4 = (({1{((-4'sd2)|(5'd0))}}+((-2'sd0)+(-2'sd1)))>({3{(5'd24)}}!=((5'd30)>(5'd4))));
  localparam signed [5:0] p5 = (((-5'sd7)+(-4'sd1))|((-3'sd3)>>(3'd4)));
  localparam [3:0] p6 = ((~&(&((5'sd10)<<<(4'd7))))?(((-4'sd6)>=(3'sd2))!==((-2'sd1)||(5'd15))):((4'd9)?(4'sd2):(3'd6)));
  localparam [4:0] p7 = (~&(~^(+(^(-(-(!(~&(+(3'd6))))))))));
  localparam [5:0] p8 = (({4{(-4'sd5)}}^(~&(2'd2)))?(~|{3{(-4'sd0)}}):{1{(^((5'd16)?(5'd2):(3'd5)))}});
  localparam signed [3:0] p9 = ({1{(((3'sd0)-(3'd2))&((4'd5)?(2'd1):(4'd10)))}}^~({4{(2'd3)}}<<<((4'sd3)==(-3'sd3))));
  localparam signed [4:0] p10 = {(3'd6),((4'd3)?(4'sd5):(-3'sd3)),((4'sd3)&(4'sd7))};
  localparam signed [5:0] p11 = ((+((5'd11)^(2'sd1)))%(-3'sd0));
  localparam [3:0] p12 = (3'd0);
  localparam [4:0] p13 = {(^(((3'sd0)?(3'd0):(3'd0))?(|(-5'sd10)):((-4'sd3)-(5'd30)))),{{((3'sd2)?(5'd30):(-2'sd0))},((3'd3)?(5'd27):(-3'sd0)),((4'd15)<<(-2'sd0))}};
  localparam [5:0] p14 = {2{((^{2{(5'd13)}})+((4'sd7)^~(-2'sd1)))}};
  localparam signed [3:0] p15 = (6'd2 * (^{(5'd19),(2'd0),(4'd14)}));
  localparam signed [4:0] p16 = (~|({1{{3{(3'd5)}}}}||((-3'sd1)-(2'd3))));
  localparam signed [5:0] p17 = ((((-3'sd1)?(5'sd5):(3'sd3))&(3'd6))>({4{(5'sd8)}}!=((5'd11)?(2'sd0):(-5'sd9))));

  assign y0 = {(+($unsigned(p3)<<(b3<=a1))),{(a1|a0),(|(a4<=p5))},{{a3,b0,b5},(p11!=a4)}};
  assign y1 = (~{3{{1{((&a0)?(p3?a1:p5):{2{b0}})}}}});
  assign y2 = (5'd0);
  assign y3 = ((b0===b5)?(p3?p7:p11):(~(p15)));
  assign y4 = ((~&(~((a0!==b1)>=(b4>b2))))===((|(a4|a1))<=(~^(^a0))));
  assign y5 = {(a0!=a1),(p5||p0),(p9^b2)};
  assign y6 = ((-2'sd0)>>(4'sd6));
  assign y7 = (|(4'd8));
  assign y8 = ((2'd2)<<<{4{(-2'sd0)}});
  assign y9 = {(~$unsigned(((-{1{p7}})))),(^(~(+{4{p6}}))),(~|{1{{(^p5),{p5,p10,p2}}}})};
  assign y10 = {1{(&$signed({3{$signed(a1)}}))}};
  assign y11 = ((6'd2 * (a2^~a0))>=(3'd0));
  assign y12 = ({(|p0),(~^p16)}?{{4{p13}},$signed(b1),$signed(p17)}:{4{a0}});
  assign y13 = ((2'd1)?{4{p1}}:{1{{4{a4}}}});
  assign y14 = $signed({2{(b1-p17)}});
  assign y15 = (b1?b2:p9);
  assign y16 = (^{2{(b3?p9:p0)}});
  assign y17 = $unsigned($unsigned($unsigned((5'd3))));
endmodule
