module expression_00648(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(3'sd2),(2'sd0)};
  localparam [4:0] p1 = ({(3'sd2)}&&((-5'sd8)+(2'sd1)));
  localparam [5:0] p2 = {2{((-4'sd0)>>(4'd3))}};
  localparam signed [3:0] p3 = (^(|(&(((5'd30)^~(-4'sd7))%(4'd0)))));
  localparam signed [4:0] p4 = {(((~|(3'd1))&{(2'd3)})<{((-2'sd0)&&(-3'sd2)),(&(3'sd3))}),(({(3'd5),(5'd21),(2'sd1)}<<((2'd2)&&(2'sd0)))&(((-2'sd0)||(-3'sd3))>>((3'd6)!=(-4'sd2))))};
  localparam signed [5:0] p5 = {{(-5'sd9)},(~(5'sd10)),((4'd4)?(2'd0):(-4'sd1))};
  localparam [3:0] p6 = (~&{{(-2'sd1),(2'd2),(2'd3)},{(3'd3),(2'd0)},{(3'sd1),(-5'sd10)}});
  localparam [4:0] p7 = {(-3'sd0),((2'd3)<<<(-2'sd0)),{(-3'sd3)}};
  localparam [5:0] p8 = (&(~|(~&((((-4'sd4)?(3'd4):(2'sd0))>((3'sd2)?(-3'sd0):(5'd15)))&(+(~(+(-4'sd3))))))));
  localparam signed [3:0] p9 = ((3'sd3)^(5'sd12));
  localparam signed [4:0] p10 = ({3{(3'd6)}}^(4'd2 * (3'd3)));
  localparam signed [5:0] p11 = (((4'sd2)?(4'd0):(5'd5))?(((-5'sd10)>>(-3'sd0))==(6'd2 * (5'd4))):(((3'd3)&(3'sd0))-((2'd0)?(4'd7):(3'd4))));
  localparam [3:0] p12 = (({(5'd30),(2'd1)}^{(2'd3),(5'd13),(2'd0)})>>>(((-4'sd3)^(2'sd1))-((2'sd1)>>>(-3'sd0))));
  localparam [4:0] p13 = (4'd5);
  localparam [5:0] p14 = ((2'd3)|(3'd0));
  localparam signed [3:0] p15 = (-(((5'd5)|(4'sd6))&((5'd24)>(-2'sd0))));
  localparam signed [4:0] p16 = {1{((3'd6)|(3'd1))}};
  localparam signed [5:0] p17 = (!{3{((2'd3)>>>(4'd9))}});

  assign y0 = (-(4'sd6));
  assign y1 = (+((b3-b0)===$unsigned(b3)));
  assign y2 = {1{(~&(((-(-{2{b4}}))!==(|(&(~|b1))))>((~|{2{a3}})>>>({2{a0}}>>(&b3)))))}};
  assign y3 = $signed($unsigned({4{(-a2)}}));
  assign y4 = {($signed((~&$unsigned((&(a0)))))?(-({p0}==(p12?a4:b5))):((-2'sd0)==(3'd3)))};
  assign y5 = $unsigned(((((b4?a5:b5)<<{4{b5}})?((~a2)^(a4?b5:p8)):{3{b2}})));
  assign y6 = ({3{p15}}-(a3===a4));
  assign y7 = (5'sd11);
  assign y8 = (-{{{{3{b2}},{p4,b5}},{3{(a3>a0)}}},((-(~$signed((~^p15))))|$unsigned({1{(a0!==b2)}}))});
  assign y9 = ({1{$signed({((p4?a0:b3)<(a4&&p12)),(p14?p10:b3)})}});
  assign y10 = $unsigned((b4^~p6));
  assign y11 = (b5<b3);
  assign y12 = ((b5!=a5)!=(3'sd1));
  assign y13 = (^((~^(^(p15?p13:p1)))?(~((&p9)%p8)):(|(~^(~|(~|p17))))));
  assign y14 = {{3{p15}},$unsigned(a0)};
  assign y15 = ({{a0}}>>(b4<=a3));
  assign y16 = (-3'sd0);
  assign y17 = {p5,p7,b0};
endmodule
