module expression_00276(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(~(!{{(4'd10)},((-2'sd0)?(4'd2):(5'd15))})),{(-{((-4'sd4)?(-2'sd0):(5'd11)),((5'd13)?(2'd1):(5'd17)),(~(2'd0))})}};
  localparam [4:0] p1 = ((-3'sd1)!==(-2'sd0));
  localparam [5:0] p2 = ({3{(-5'sd4)}}>>>{1{(-5'sd9)}});
  localparam signed [3:0] p3 = {1{((-4'sd4)!=(2'd2))}};
  localparam signed [4:0] p4 = {(|{(3'd6),(^((-3'sd3)!=(-4'sd2)))})};
  localparam signed [5:0] p5 = ((((3'sd1)>=(3'd4))===(|(-(-2'sd0))))!==(+(^(!(2'd3)))));
  localparam [3:0] p6 = ({3{(5'sd3)}}!=={3{(2'sd0)}});
  localparam [4:0] p7 = (((-4'sd7)+(2'd2))|((4'sd7)?(5'sd1):(4'd7)));
  localparam [5:0] p8 = (5'd5);
  localparam signed [3:0] p9 = (((3'd5)^~(-5'sd1))*((5'sd1)==(5'sd2)));
  localparam signed [4:0] p10 = {(((6'd2 * (5'd15))?(-5'sd0):{1{(3'd0)}})&({(5'd10),(4'sd1),(3'sd1)}^((2'sd0)?(5'sd7):(4'sd3))))};
  localparam signed [5:0] p11 = ((!(-3'sd3))===((2'd3)>>>(2'sd0)));
  localparam [3:0] p12 = {{((5'sd13)^(4'd13)),{(2'd3)},((2'd3)^(3'sd3))},{((5'sd3)?(5'd28):(4'd5)),((4'sd6)?(3'd0):(4'sd4))}};
  localparam [4:0] p13 = ((2'd2)!=={2{{3{(3'd1)}}}});
  localparam [5:0] p14 = {3{{((5'sd3)?(4'sd7):(5'd27))}}};
  localparam signed [3:0] p15 = (~|(~&(|((-4'sd0)%(2'sd0)))));
  localparam signed [4:0] p16 = (((5'd11)<=(4'd1))?((3'sd3)^~(3'd3)):{4{(2'd0)}});
  localparam signed [5:0] p17 = (5'sd6);

  assign y0 = (-4'sd2);
  assign y1 = ((b1==p11)+(~&(~a4)));
  assign y2 = (((-(4'd13))/p3)!=(-4'sd5));
  assign y3 = {2{(3'd3)}};
  assign y4 = ({1{(!(|(+{1{{1{$unsigned($unsigned(p11))}}}})))}});
  assign y5 = (((p12-p10)?(b0|p10):(p15<p2))?(!((p10?a2:p2)?(p14!=p7):(p15?p3:p11))):((p13^p14)*(4'd2 * p12)));
  assign y6 = (5'd26);
  assign y7 = {4{(^{2{b0}})}};
  assign y8 = ((p4>=p11)%a0);
  assign y9 = {((~^(p16&p16))?($signed(p5)):(a0===b5)),(-(((p13&p14))<<(!(~p11))))};
  assign y10 = (p15>a3);
  assign y11 = ({{1{(b3&a4)}},{b1,b2},{{1{p2}}}}&&(($unsigned({4{a2}}))<<({a3}>>>(b3<b3))));
  assign y12 = ((3'd3)>>>(b1^p2));
  assign y13 = (+(^(~^(~^(-{(&(+(b1<<<b5))),((!a1)!==(^a1)),{(a2<a0)}})))));
  assign y14 = ({3{a0}}-{2{b1}});
  assign y15 = (p4);
  assign y16 = $signed(({4{{(p3<<<a5)}}}|$unsigned(({4{a3}}<<((a0&&b0)!==(a4+a0))))));
  assign y17 = (|(^(-(&(+(-{2{$signed($unsigned((~|(!(!p11)))))}}))))));
endmodule
