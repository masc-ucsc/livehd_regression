module expression_00438(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-3'sd3);
  localparam [4:0] p1 = ((((-3'sd2)?(-5'sd4):(-4'sd3))<((-2'sd0)?(2'sd1):(2'd2)))!=(((3'd0)+(5'd2))?((4'd7)>>(5'd12)):((4'd3)!=(5'd28))));
  localparam [5:0] p2 = (3'd6);
  localparam signed [3:0] p3 = (({1{(^(3'd5))}}==((5'sd11)?(5'sd14):(-2'sd0)))<<{2{(+(+(-4'sd3)))}});
  localparam signed [4:0] p4 = (|((((4'd10)||(5'd30))+(~((2'd3)!=(5'd4))))^(-(((4'd9)>>>(5'd23))>>((-5'sd10)-(4'd7))))));
  localparam signed [5:0] p5 = (((2'd1)?(4'd12):(3'd2))/(2'd0));
  localparam [3:0] p6 = ({3{((5'd12)!=(4'sd7))}}<=(((3'd4)-(-3'sd3))&&{1{(3'sd0)}}));
  localparam [4:0] p7 = ({((2'd3)-(5'd12)),((4'd0)>>(3'sd3))}==((5'd2 * (3'd6))&{(-2'sd0),(3'd6)}));
  localparam [5:0] p8 = {4{((2'sd1)&&(3'd1))}};
  localparam signed [3:0] p9 = (~(5'd8));
  localparam signed [4:0] p10 = (~&(&(3'd2)));
  localparam signed [5:0] p11 = ((((3'sd2)?(4'd9):(2'd2))?((3'd4)?(5'd27):(-2'sd0)):{1{(2'sd0)}})?(!(~|((5'd6)?(-4'sd3):(3'd2)))):{2{((3'd3)?(-5'sd1):(2'd0))}});
  localparam [3:0] p12 = {((2'sd1)>={(5'sd8),(2'd1)}),{{3{(3'sd1)}}},({(3'sd3),(-2'sd0),(2'd1)}^{(2'd1)})};
  localparam [4:0] p13 = ((((5'd12)-(2'sd1))>={1{(4'sd4)}})>((~&(5'd15))<<((3'd7)&(4'sd5))));
  localparam [5:0] p14 = {{{(2'sd1),(5'd4),{(4'd0),(3'd7),(3'sd1)}}},{{(-4'sd2),(2'd2),(-3'sd1)}}};
  localparam signed [3:0] p15 = (-(3'd6));
  localparam signed [4:0] p16 = ((2'd1)?(3'd2):(-4'sd5));
  localparam signed [5:0] p17 = (5'sd6);

  assign y0 = (a1<b4);
  assign y1 = ((~((-4'sd7)>>(a3-a2)))===(-2'sd0));
  assign y2 = {{2{a2}},(a5<=b1)};
  assign y3 = (2'd1);
  assign y4 = (($signed(((-2'sd1)-{{a3,a0,a3}})))<$signed({((p9>=a3)>>>(p15^~p10))}));
  assign y5 = (~(|((~|(|(a5+p4)))!={1{(p2||p1)}})));
  assign y6 = (((&(a0?p3:b2))?(3'sd1):(4'sd6))==((a3<<<a5)?(+(b2<=a0)):(b5+a2)));
  assign y7 = ({4{(5'd2 * b1)}}<<<((~&{b0,a0,b2})<{4{p17}}));
  assign y8 = ({(5'd13),$signed(b3),(3'sd2)}==={(~(~&(|$unsigned(a2))))});
  assign y9 = ({p5,b0}>>>{4{p3}});
  assign y10 = (+(4'sd6));
  assign y11 = $unsigned(((~($signed(p12)?(a5>>>b5):(6'd2 * p2)))<<<(|((6'd2 * p14)<{a2,b2}))));
  assign y12 = ((~(^(+((p7?p12:p1)>(p13<=b5)))))?(~^((p5||p2)|(^(p7<p16)))):((p16?p9:p14)!=(~&(&p11))));
  assign y13 = (6'd2 * (~{2{p6}}));
  assign y14 = ((5'sd14)?(p4?p13:p3):{p1});
  assign y15 = (4'sd2);
  assign y16 = (({p2}>>>{4{p2}})>{3{{p4,p16,p17}}});
  assign y17 = (((~|(~a0)))?(&(p2?p4:b1)):{$unsigned(p13),(-p13)});
endmodule
