module expression_00681(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((4'sd4)?(3'd3):(2'd0))<<(3'sd0));
  localparam [4:0] p1 = (((2'd3)?(-3'sd2):(-4'sd1))?((4'd0)?(2'sd0):(5'sd10)):((2'sd1)?(3'sd2):(3'd0)));
  localparam [5:0] p2 = (((5'd5)&(-5'sd5))<=((-2'sd0)?(4'd7):(5'd18)));
  localparam signed [3:0] p3 = ((5'sd3)?(2'd1):(2'sd1));
  localparam signed [4:0] p4 = (~&{2{{3{((-2'sd0)-(4'd1))}}}});
  localparam signed [5:0] p5 = {2{{3{(5'd22)}}}};
  localparam [3:0] p6 = (((5'sd10)?(4'sd4):(5'd8))?{1{{(3'd2),(2'd3)}}}:{(2'd0),(2'sd1),(5'd8)});
  localparam [4:0] p7 = {3{(((4'd3)^~(2'd1))||((-2'sd1)>>(2'd1)))}};
  localparam [5:0] p8 = ((2'd3)>>>(5'd26));
  localparam signed [3:0] p9 = (|(~^(~|((-(5'd12))=={(5'd16),(2'd0),(3'd1)}))));
  localparam signed [4:0] p10 = (~^(((2'd0)?(-5'sd10):(-5'sd7))<={2{(3'd7)}}));
  localparam signed [5:0] p11 = {4{(~^{1{{1{(2'd1)}}}})}};
  localparam [3:0] p12 = {4{{1{(^((4'd3)?(5'd7):(4'd10)))}}}};
  localparam [4:0] p13 = ((4'd2)<<<(3'd4));
  localparam [5:0] p14 = (2'd3);
  localparam signed [3:0] p15 = {2{((|(-3'sd3))===(~&(4'sd0)))}};
  localparam signed [4:0] p16 = ((5'd2 * (5'd3))<<<((4'd5)!==(-5'sd2)));
  localparam signed [5:0] p17 = (~&(((4'd13)==(3'd3))>>{(2'sd0),(-3'sd1)}));

  assign y0 = $unsigned(({4{(3'd3)}}+(2'd2)));
  assign y1 = (+(^(&(~|(~(+(~a5)))))));
  assign y2 = (~^{4{(b4?b3:p10)}});
  assign y3 = (~|{2{({{{b0,a0}}}==={(-3'sd3)})}});
  assign y4 = (((p0>>>a5)?(p3-p10):(4'd3))?((a2?p13:p13)?(4'd14):{4{a2}}):((b0>a4)!==(b4==a2)));
  assign y5 = {1{{(a2+b0),(b3&&p9),(p4?a2:p11)}}};
  assign y6 = ({(~&(&(p7!=p4))),$unsigned({(&p7)})}<<<(((&a5)||{p3})>>({p4}||$signed(p6))));
  assign y7 = ((&((p5?p17:a5)?(a1&b0):(~|(3'd3))))>>>{1{((-4'sd0)-(!(a1<a0)))}});
  assign y8 = ($signed(p1)?(p12?p7:p11):{3{p1}});
  assign y9 = ({(p15^~p14),{4{p9}},{4{p5}}}||{{3{p8}},{p3,p11},{p8,p2}});
  assign y10 = (-{1{(((a5||b4)<{2{a4}})&&((!(p10<=p13))!=(b1===a5)))}});
  assign y11 = {1{(a2||b1)}};
  assign y12 = $signed(({1{(-5'sd11)}}));
  assign y13 = {((3'sd1)<=(^(b4<<p15))),(~|(3'd3)),((a2^p10)!=(2'd3))};
  assign y14 = $signed(((~&{(p12^p10),{p16,p5,p7}})));
  assign y15 = (3'sd1);
  assign y16 = (&(p9%p2));
  assign y17 = (|((~p4)?(a0|p16):(&a2)));
endmodule
