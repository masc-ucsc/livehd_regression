module expression_00722(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((((4'd5)>>(-4'sd7))==={(-3'sd0),(4'd7)})!=={((-3'sd2)&(3'd3)),((3'd5)^~(4'sd7))});
  localparam [4:0] p1 = {2{(2'd0)}};
  localparam [5:0] p2 = ((4'd14)|(-3'sd1));
  localparam signed [3:0] p3 = ((5'd2 * ((3'd4)|(5'd19)))>((((4'sd4)&&(5'sd8))-((-3'sd1)^~(3'd4)))<(((5'd1)|(3'sd0))||(5'd2 * (5'd21)))));
  localparam signed [4:0] p4 = (((+(2'd1))?{4{(5'd21)}}:((-5'sd4)&&(-3'sd0)))>=({3{(3'd5)}}&&(~|(!(4'sd4)))));
  localparam signed [5:0] p5 = (3'sd2);
  localparam [3:0] p6 = (4'd2 * (~^(5'd12)));
  localparam [4:0] p7 = (!((|((~(5'sd6))<(&(5'sd2))))<((+(3'd0))>>((3'd0)!=(-3'sd2)))));
  localparam [5:0] p8 = (((5'sd8)&&(3'd2))*((2'd3)>(5'd28)));
  localparam signed [3:0] p9 = {{2{(3'sd2)}},{4{(3'sd2)}}};
  localparam signed [4:0] p10 = (&{((-5'sd12)<=(3'sd0)),((3'd6)>=(3'sd0)),{((3'd3)<=(3'd5))}});
  localparam signed [5:0] p11 = (((2'd1)>(2'd3))|{(4'sd4)});
  localparam [3:0] p12 = (~|({(4'sd0),(5'd27)}^(~&(~&(2'sd0)))));
  localparam [4:0] p13 = (((^(2'd1))&&{(-2'sd0),(-3'sd3)})?((2'd0)?(2'd2):(5'd9)):((|(5'd30))&&(&(2'd2))));
  localparam [5:0] p14 = (((4'd14)<<(-2'sd0))&((-5'sd13)?(2'd2):(3'd0)));
  localparam signed [3:0] p15 = {2{{1{(5'sd15)}}}};
  localparam signed [4:0] p16 = (((3'd0)+(-2'sd0))^((5'd8)!==(4'sd5)));
  localparam signed [5:0] p17 = (~&({{(2'sd1),(4'sd2)},((2'd2)<(4'sd2)),((5'sd9)!==(2'sd0))}!==(((4'sd3)>=(-3'sd3))+(^(+(4'd9))))));

  assign y0 = {{{a3,a1},(!b1),$signed(b5)},$signed($signed((|(|{p2,p14,p15}))))};
  assign y1 = {3{{2{(~^{b5})}}}};
  assign y2 = (&(4'sd0));
  assign y3 = {4{(a3>>p9)}};
  assign y4 = ((p5>>>b3)>(a3|p1));
  assign y5 = (5'd2 * (b0^p1));
  assign y6 = (^((+(5'd22))>=(b4-b4)));
  assign y7 = ((2'd2)||{(2'd2)});
  assign y8 = ((6'd2 * (b2>p1))?(-((&a1)!=={1{b1}})):(+{4{p0}}));
  assign y9 = ({$unsigned({3{b1}}),$signed((~p5)),(&(p14))});
  assign y10 = {(~{(+(3'd4))})};
  assign y11 = {({(~p5)}^(p14>b0))};
  assign y12 = (~|(((b3||a4)^~(a2<=a3))>>(~|((~(b1===a2))===(b2<a5)))));
  assign y13 = (~^((b3===a5)||(b2|b1)));
  assign y14 = (4'd5);
  assign y15 = ((((-b5)>(a4==b3))&&((-5'sd2)>>(+a3)))===((-(a3<=b2))!==(|(|(b0!=a3)))));
  assign y16 = ((p13?p6:p7)?(~|$signed((&p0))):(&(~(a0!=p17))));
  assign y17 = ((a4^~b1)?(3'sd1):(b2?b5:b0));
endmodule
