module expression_00435(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((3'd1)?(((2'sd0)?(-4'sd1):(4'd11))==((4'd2)?(4'd8):(4'd10))):(3'd0));
  localparam [4:0] p1 = {3{{4{(5'd28)}}}};
  localparam [5:0] p2 = ({(4'd2),(4'sd1),(5'd12)}^~((5'd31)<<<(5'sd15)));
  localparam signed [3:0] p3 = (((3'd0)<(3'sd0))?((-3'sd1)?(-3'sd0):(2'd3)):((3'd6)<(5'sd10)));
  localparam signed [4:0] p4 = (~^{(|((!(2'd1))==(|(5'd24))))});
  localparam signed [5:0] p5 = ((((2'd0)?(-2'sd0):(-5'sd15))+(&{((5'd15)<=(5'sd1))}))>((-((-4'sd6)?(4'sd5):(-3'sd2)))<<(-((5'sd2)>>>(-2'sd0)))));
  localparam [3:0] p6 = {1{({3{{1{(5'd5)}}}}-{2{{1{(-4'sd3)}}}})}};
  localparam [4:0] p7 = (((^{(3'd6),(3'd5)})<<{4{(2'd3)}})&({(5'sd9),(2'd1)}>>((5'sd12)>=(5'd10))));
  localparam [5:0] p8 = (6'd2 * ((4'd2)<=(2'd2)));
  localparam signed [3:0] p9 = ({4{(2'sd0)}}=={1{((-(-4'sd3))==(3'd4))}});
  localparam signed [4:0] p10 = {(^((2'd0)?(2'sd0):(2'd3))),(((-2'sd0)?(4'd14):(4'd1))>>>(&(4'd0))),{((4'd0)?(2'd1):(-4'sd7)),((3'd1)?(-3'sd3):(2'sd0))}};
  localparam signed [5:0] p11 = {{{{({(-2'sd0)}+((3'd0)||(2'sd1)))}}}};
  localparam [3:0] p12 = (((3'd7)?(4'sd7):(-3'sd3))?{4{(5'd3)}}:{4{(-2'sd1)}});
  localparam [4:0] p13 = ((-3'sd3)!=(4'd12));
  localparam [5:0] p14 = (+{4{((~(-3'sd3))||(&(-5'sd8)))}});
  localparam signed [3:0] p15 = (3'd6);
  localparam signed [4:0] p16 = (((-4'sd6)?(2'd0):(4'sd1))?((5'sd15)?(4'd14):(5'd27)):((5'sd15)==(4'd4)));
  localparam signed [5:0] p17 = (((4'd6)+(3'sd1))<<((2'd3)<=(-2'sd0)));

  assign y0 = (5'd9);
  assign y1 = (&(((~|(p3<<a5))%a2)?(~^((p15?p0:b2)/a3)):((a1==a3)===(b1|a1))));
  assign y2 = ({{a3,b3,a3},(b3||p15),{4{b0}}}^~{(((p15))),{4{b1}}});
  assign y3 = (~&(-(((!(~|(~|b4)))<=((|a3)&&(+b2)))&(((a5!=p11)^~(+a4))<<<(&(a1^a0))))));
  assign y4 = ((p6?p16:p2)%p1);
  assign y5 = (((a2?a3:a0)^~(b2?b0:b3))?((b3<<b1)&&(b3?b2:b3)):(6'd2 * (b1<=a2)));
  assign y6 = (({b3,p2})<{(&b5)});
  assign y7 = (-3'sd3);
  assign y8 = (~&(~|b3));
  assign y9 = (((4'sd1)?(b2^~a1):(-5'sd14))?((a4^p13)+(5'd5)):((a2<<<b2)==(5'sd9)));
  assign y10 = (~(~^(~^{4{(-(5'sd11))}})));
  assign y11 = $signed((|{(p7>p12),{$unsigned(p17)},{p4,p13}}));
  assign y12 = ((((b1^a5)||(a5<<a3))<<<((a5<b3)<<(b4&a1)))^~(((p3/b1)/p14)|((a4>a0)>(p16==p3))));
  assign y13 = ((~|((p9>>p17)<<{3{a2}}))<=((-(b0^p3))||({3{p11}}>>(b5!==a4))));
  assign y14 = (~^(~^(~|(((~&(4'd2 * p8))>>((b1===a1)>>(~^a4)))<<(((p10^~p7)<=(|p0))<=((|a0)===(b4^~a1)))))));
  assign y15 = ((|((^(a5>>a4))|(b4===b5)))^~(+((p3||b1)^(b2/a1))));
  assign y16 = {1{((~({2{(~^{3{a5}})}}|(((~|p1)|{3{p0}})))))}};
  assign y17 = (~^((~^((~p5)?(^p5):(~|b5)))<<<{2{(+{2{b5}})}}));
endmodule
