module expression_00253(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (&(({3{(-3'sd3)}}?(~(-5'sd6)):(~|(5'sd10)))>(4'd2 * (-{1{(3'd5)}}))));
  localparam [4:0] p1 = (|(-(~&(&({1{{3{(-2'sd1)}}}}?{(4'd3),(5'sd12),(5'd19)}:{1{(~|(2'd1))}})))));
  localparam [5:0] p2 = {(~&{((-5'sd2)?(2'd3):(-4'sd3)),{2{(5'd6)}}})};
  localparam signed [3:0] p3 = (^(~^((&(4'sd0))<=(|(3'd3)))));
  localparam signed [4:0] p4 = (-{2{(4'd8)}});
  localparam signed [5:0] p5 = ({(3'sd1),(5'd6)}<((3'sd1)<=(2'sd1)));
  localparam [3:0] p6 = (~{{(-(-2'sd0)),{(3'sd1),(-5'sd15)}},(((-4'sd3)^(2'd3))<=(!(2'd1)))});
  localparam [4:0] p7 = (!(&(&(-4'sd7))));
  localparam [5:0] p8 = {({(-4'sd2),(-5'sd4),(4'd13)}!=((-3'sd3)&(5'd26))),{2{((5'd4)<=(5'd9))}}};
  localparam signed [3:0] p9 = {3{{1{(-5'sd6)}}}};
  localparam signed [4:0] p10 = (~^(&(-3'sd2)));
  localparam signed [5:0] p11 = {1{{3{({1{(-4'sd0)}}-{2{(4'd4)}})}}}};
  localparam [3:0] p12 = (4'sd3);
  localparam [4:0] p13 = (!((((5'd26)||(-5'sd6))^~(|(-5'sd9)))^~(|{(^(~(-2'sd1)))})));
  localparam [5:0] p14 = ((3'sd0)?(-2'sd0):(4'sd2));
  localparam signed [3:0] p15 = (6'd2 * ((5'd24)?(3'd4):(3'd5)));
  localparam signed [4:0] p16 = {{(&(~|((5'd31)>>>(4'sd1)))),(|(^((3'd5)^(3'd6))))}};
  localparam signed [5:0] p17 = ((6'd2 * (2'd2))?((4'd6)&(4'sd0)):((5'd12)?(-2'sd0):(3'sd3)));

  assign y0 = (~&(&((^($signed(b5)^~(b5)))&&(~|((&a0)|(a3^a1))))));
  assign y1 = {4{(p16|p4)}};
  assign y2 = (-((-(^(5'd2)))?(5'd12):{3{(b3?p2:p0)}}));
  assign y3 = ((a4&p14)+$unsigned((&b1)));
  assign y4 = (({1{(~^(2'sd1))}}^~(~|(b1>>>b4)))<=((5'd16)-((2'sd1)^~(p7?p8:b3))));
  assign y5 = ((+(!((|a1)?(a0?b2:p3):(b0-a3))))-{({b1}?(b1?a2:b0):(-a0))});
  assign y6 = $signed((~|$unsigned(((~&$unsigned(b0))?(|$unsigned(p6)):(p1>>>a3)))));
  assign y7 = (|(&(~&p12)));
  assign y8 = (3'd1);
  assign y9 = {1{{2{(~(~^(~(-(|b0)))))}}}};
  assign y10 = (((~p16)?(a3>a4):(a3?a5:p6))^((~(a1<a5))^(~^(+a4))));
  assign y11 = (~&{1{(~|b1)}});
  assign y12 = (a0<<<b4);
  assign y13 = (a3===b4);
  assign y14 = ({4{(a0?b2:a2)}}<=((b1?b1:a1)==={2{a3}}));
  assign y15 = (~^((p8==p15)|{p1}));
  assign y16 = (((4'd0))<=($signed({a2,a2,p11})+{p9,p13,p1}));
  assign y17 = (((b2?a3:a5)*(a2!=a3))&&(~^(~|(4'sd0))));
endmodule
