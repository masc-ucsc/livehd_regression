module expression_00882(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (!(-3'sd1));
  localparam [4:0] p1 = ((-2'sd0)?(2'd0):(4'd8));
  localparam [5:0] p2 = (&(~&(+(5'sd5))));
  localparam signed [3:0] p3 = (~|(!(^(~&(~|(5'd18))))));
  localparam signed [4:0] p4 = (!(((4'sd2)>(-4'sd4))*(~^(~&(-2'sd0)))));
  localparam signed [5:0] p5 = {((4'd8)?(-2'sd0):(4'd7))};
  localparam [3:0] p6 = ((~^(5'sd6))<=(~&(3'd4)));
  localparam [4:0] p7 = (((4'd2 * (4'd7))/(4'd1))>>(((4'sd1)+(4'd12))^~((2'd0)+(5'd13))));
  localparam [5:0] p8 = ((-(3'd6))?((-4'sd1)?(5'd6):(3'd7)):(|(4'sd7)));
  localparam signed [3:0] p9 = (|(((5'sd13)?(3'sd0):(5'sd14))?((3'sd0)?(-4'sd3):(3'd7)):((2'd0)?(2'sd0):(-4'sd4))));
  localparam signed [4:0] p10 = {1{{4{(4'd12)}}}};
  localparam signed [5:0] p11 = (-2'sd0);
  localparam [3:0] p12 = (+(5'd2 * {3{(4'd1)}}));
  localparam [4:0] p13 = (((4'sd3)<<(5'sd14))?((-5'sd8)?(3'sd3):(3'd0)):(4'd2 * (5'd18)));
  localparam [5:0] p14 = (&{2{(|{4{(2'd2)}})}});
  localparam signed [3:0] p15 = (|{3{(3'd0)}});
  localparam signed [4:0] p16 = (~|((!(3'd0))<<<(3'sd1)));
  localparam signed [5:0] p17 = {(~{(5'd22),(4'sd4),(4'sd7)}),{((-4'sd2)?(3'd1):(2'd0))},(~&(-((5'd18)==(-5'sd5))))};

  assign y0 = (((+(a5-a0))?(p7<<<p9):(a1^~b5))<<{(((~^b3)|{b1,p0})<=(~(b3!==a1)))});
  assign y1 = (-a5);
  assign y2 = {((p7>>p15)==(a5?p2:p2))};
  assign y3 = (((3'sd1)||(p1/p16))|(5'sd10));
  assign y4 = $signed((&((3'sd1)|((-5'sd0)/a5))));
  assign y5 = $unsigned($signed($unsigned((($signed($unsigned(($signed($unsigned(($signed($signed(a4)))))))))))));
  assign y6 = (&(!b3));
  assign y7 = (+((~|(a0?a5:a3))!==(b0?b0:a2)));
  assign y8 = {(-5'sd14),$unsigned($unsigned(((b1-a1)===(-b0)))),((b0!=a3)!=(b2||p11))};
  assign y9 = (~^(|p16));
  assign y10 = (2'd1);
  assign y11 = (3'd0);
  assign y12 = $unsigned((~&a1));
  assign y13 = (5'sd0);
  assign y14 = ((~^((b0?a0:a0)&&(-a1)))-(-(|(6'd2 * b2))));
  assign y15 = ({{1{a5}}}?(5'd2):{(p17?p6:p16)});
  assign y16 = (+(((2'sd0)^~(4'd2 * p6))<=(~{(|(p7))})));
  assign y17 = {(&{2{(^({2{a5}}>={a2,a2}))}})};
endmodule
