module expression_00724(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~^(2'sd0));
  localparam [4:0] p1 = (~{((!((4'sd0)?(-4'sd1):(-4'sd2)))&(((5'd23)?(5'd2):(4'd11))?((-5'sd1)|(-5'sd0)):((-3'sd2)-(3'sd3))))});
  localparam [5:0] p2 = ({{3{(-2'sd0)}},{(2'sd1),(-3'sd2),(-4'sd1)}}<<({4{(-2'sd0)}}>>>((3'd5)?(4'd5):(2'd2))));
  localparam signed [3:0] p3 = (((3'sd2)|(4'd11))^~(-(-5'sd7)));
  localparam signed [4:0] p4 = (~(-2'sd0));
  localparam signed [5:0] p5 = ({(-4'sd3),(5'd24),(2'sd1)}>({(4'd11),(5'sd11)}&{(2'd2),(3'sd0)}));
  localparam [3:0] p6 = {(((5'sd4)>>>(-4'sd3))<=((4'd2)<<(4'd11))),(^(4'd2 * ((2'd0)>>(3'd2))))};
  localparam [4:0] p7 = {(4'sd5),{{(-3'sd3),(2'd1)},((5'd30)&&(-3'sd3))}};
  localparam [5:0] p8 = (~((~((5'sd13)===(2'd1)))?(-(-4'sd4)):(-5'sd4)));
  localparam signed [3:0] p9 = {(~(4'd10)),((3'd1)!=(4'sd7)),((2'd3)^(5'd14))};
  localparam signed [4:0] p10 = {(-4'sd0),(((2'd2)|(3'sd2))|{(-2'sd0),(-4'sd7)}),(3'd4)};
  localparam signed [5:0] p11 = (~&(~({((~^(3'd7))!=((4'd3)>>>(3'd2)))}-({(5'd21),(4'd10),(-2'sd1)}&((3'd7)^(4'd2))))));
  localparam [3:0] p12 = ({1{{((2'd3)>(-3'sd0))}}}>=(5'd10));
  localparam [4:0] p13 = ((-2'sd0)!==(5'd4));
  localparam [5:0] p14 = (|(^(((5'd29)<=(2'd1))?((5'sd4)>>>(3'd4)):((2'd3)<=(5'd5)))));
  localparam signed [3:0] p15 = {{(~&(5'sd9)),(+(-3'sd1)),(+(3'd2))},(!{{(4'd12)},(~^(4'sd6))})};
  localparam signed [4:0] p16 = (&(-((4'd10)-(-4'sd4))));
  localparam signed [5:0] p17 = (6'd2 * ((3'd2)<=(2'd0)));

  assign y0 = (+((-(&(~^(a4>>a4))))&(~&((!a1)|(-a1)))));
  assign y1 = ({3{{2{b5}}}}||(-$signed({{4{(p0||p11)}}})));
  assign y2 = (-3'sd2);
  assign y3 = {3{(~&{1{$unsigned({2{a4}})}})}};
  assign y4 = ((b4+p16)<<(p11/p1));
  assign y5 = (-4'sd0);
  assign y6 = ({3{a2}}^(b3>>a1));
  assign y7 = ((p1?p16:b5)?{1{(3'd0)}}:(~^(p13?p14:p14)));
  assign y8 = (2'd2);
  assign y9 = {2{({(4'd10)}>=(b4||b4))}};
  assign y10 = {((~{b3})===(a2<=b2)),(5'd27),(+(-(&(|{p17,b5,b2}))))};
  assign y11 = {((2'd3)+(a0-p2)),{(2'd1),(5'sd13)},((a1?p4:a1)-(~p8))};
  assign y12 = {(~^(^(2'd3))),{(~(~&(3'sd3)))}};
  assign y13 = (p16>>>p0);
  assign y14 = {p11,b5};
  assign y15 = ((2'sd1)&&{2{((-3'sd2)<<(b1?b0:b1))}});
  assign y16 = {3{(a2^~p1)}};
  assign y17 = (2'sd0);
endmodule
