module expression_00331(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(-5'sd12),(-5'sd3)};
  localparam [4:0] p1 = (^(^(-(~|(~^((-(|(^(5'd10))))<(-(~{2{(4'd7)}}))))))));
  localparam [5:0] p2 = ((((4'sd7)>(-4'sd1))!=((3'sd0)<=(-4'sd6)))&&(((3'd5)%(5'd10))!=((-3'sd0)|(-5'sd9))));
  localparam signed [3:0] p3 = ((((2'd1)&&(4'd7))-(5'sd3))<<(!(2'd0)));
  localparam signed [4:0] p4 = (!((~&((-4'sd6)>(5'sd11)))>=((5'sd11)>(2'd0))));
  localparam signed [5:0] p5 = (4'd2);
  localparam [3:0] p6 = ((((4'sd6)==(-5'sd12))>>>((5'd17)<(-3'sd1)))+(((5'd1)<<<(-2'sd1))-((-4'sd0)+(2'sd1))));
  localparam [4:0] p7 = (3'd3);
  localparam [5:0] p8 = ({4{(4'd7)}}?{2{((5'sd13)?(5'sd15):(-5'sd4))}}:{4{(-4'sd6)}});
  localparam signed [3:0] p9 = ({(4'd8),(5'd3),(-2'sd1)}-((3'd1)&&(-4'sd0)));
  localparam signed [4:0] p10 = (-((((-5'sd8)|(3'sd1))&&{(5'sd5)})|{((3'd2)&(3'd4)),{2{(-2'sd1)}}}));
  localparam signed [5:0] p11 = ((2'sd1)-((5'sd15)==(2'sd0)));
  localparam [3:0] p12 = ((((4'd10)!=(-4'sd0))&((5'd6)+(2'd0)))-({2{(-5'sd14)}}>>>((5'sd11)==(3'd5))));
  localparam [4:0] p13 = (((2'd2)&(2'd1))<=(~|(3'd6)));
  localparam [5:0] p14 = (3'sd3);
  localparam signed [3:0] p15 = (((3'd6)<<<(5'd15))?((-3'sd2)^(5'sd9)):(+(5'd1)));
  localparam signed [4:0] p16 = (~^(~|(~(((4'd1)?(-2'sd1):(3'd2))?((3'sd0)>>>(5'd15)):((2'sd0)<<<(3'sd0))))));
  localparam signed [5:0] p17 = ((^(~^(4'd9)))%(-2'sd1));

  assign y0 = (((p10<=p1)-(-(p11+p5)))||((!(p16!=p16))<=(p6||p17)));
  assign y1 = (!((~^(~&(&(+(p5?b4:a4)))))?({p9}?{p14,b1}:(b1?b4:p0)):({a2,p12}&&(|(&p17)))));
  assign y2 = $unsigned((~|(-2'sd0)));
  assign y3 = (~p2);
  assign y4 = (~a3);
  assign y5 = (+$signed((|(b1!==b3))));
  assign y6 = {2{((a1?p6:a3)?(p11^b0):(-(+p16)))}};
  assign y7 = $unsigned(p0);
  assign y8 = ((!{3{p2}})?{3{p15}}:{3{a3}});
  assign y9 = {({(a4+b4),{a3},(a2^~a4)}!==({b4}==={a0}))};
  assign y10 = (((b1)/p12)&&($unsigned(a5)!==(b2>>>b5)));
  assign y11 = ((((b4&a0)?{4{b3}}:(b5?b4:a0)))===({4{a3}}|((+(~^{4{a4}})))));
  assign y12 = (!(((|(^p9))?(p13||p15):{p3,p4,p17})>({(p13?p11:p11),(p13?p10:p14)}<((p14?p10:p0)&{p9}))));
  assign y13 = ({$unsigned(b1)}&(b4||p0));
  assign y14 = (-2'sd0);
  assign y15 = {(^(+(&p5))),(5'd2 * (p12<=a0)),((p12!=b0)!=(a3-b2))};
  assign y16 = (p11>>p14);
  assign y17 = ({b3,a2}?(a2<<<b0):(3'sd0));
endmodule
