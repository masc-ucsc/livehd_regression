module expression_00905(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd23)-(4'd12));
  localparam [4:0] p1 = (((-3'sd3)?(3'd4):(4'd10))?((-5'sd8)?(-5'sd2):(4'sd4)):((^(-3'sd2))===((2'd3)?(4'd0):(2'd2))));
  localparam [5:0] p2 = {2{{2{{1{{3{(3'sd3)}}}}}}}};
  localparam signed [3:0] p3 = {({4{(-5'sd7)}}===((2'sd1)!=(-3'sd3))),((~(2'sd0))>>((4'sd7)>>(-3'sd0))),(((-4'sd0)<<(4'd7))^~{(5'd0),(3'd6),(3'sd2)})};
  localparam signed [4:0] p4 = ((4'd2 * (2'd1))?((2'd2)-(-3'sd3)):((-4'sd0)?(5'sd0):(4'd10)));
  localparam signed [5:0] p5 = (4'd2 * {1{(~|(4'd5))}});
  localparam [3:0] p6 = (((2'd2)?(2'd2):(5'd24))^~((-3'sd1)?(4'sd6):(2'sd0)));
  localparam [4:0] p7 = ((-4'sd3)+{4{(2'sd1)}});
  localparam [5:0] p8 = ((-((-2'sd0)?(5'sd15):(2'd1)))&(2'sd1));
  localparam signed [3:0] p9 = {{(2'd1),(2'd3),(5'd26)}};
  localparam signed [4:0] p10 = {(^(+(+{(5'sd13),(2'd0)}))),{(^(2'd0)),(^(5'd8))}};
  localparam signed [5:0] p11 = (((-4'sd3)|(-5'sd15))?(-((3'd0)==(4'sd5))):((3'd2)>>(5'd5)));
  localparam [3:0] p12 = (-(~^((-(-(5'd7)))>>>(|{4{(2'd3)}}))));
  localparam [4:0] p13 = (~((^(~^{4{(-3'sd3)}}))>={{(3'd3),(5'd10)}}));
  localparam [5:0] p14 = (5'd11);
  localparam signed [3:0] p15 = ({4{(5'd19)}}?((5'sd6)|(2'sd0)):{(-4'sd2),(4'd0),(-3'sd3)});
  localparam signed [4:0] p16 = ((|(~(~(2'd3))))^(((3'd0)?(2'd0):(-2'sd1))|((2'sd0)?(5'sd14):(2'd0))));
  localparam signed [5:0] p17 = ({1{((4'd14)?(4'd3):(5'sd4))}}===((5'sd1)?(-3'sd3):(-4'sd0)));

  assign y0 = (4'd6);
  assign y1 = (5'sd8);
  assign y2 = $unsigned($signed($unsigned(((((($unsigned($unsigned(((b4))))))==$signed(($unsigned(($unsigned(a4)*(a4<<a4)))))))))));
  assign y3 = (~(2'sd0));
  assign y4 = {{((-{a4,p2,a1})>>(a5>b0)),({(~^p0)}<<(a2>>b2)),((^(a3>>>b4))==={1{(a0^b5)}})}};
  assign y5 = ((~&(b0?a2:b3))*(~|(b0?a5:b0)));
  assign y6 = ((a5>=p13)!={a2,b2,a1});
  assign y7 = {(a4+b0),(b4!=b1),(b1^b2)};
  assign y8 = $signed((!(-{3{{1{(&{{{p13,p6}}})}}}})));
  assign y9 = {4{a2}};
  assign y10 = (a3===a5);
  assign y11 = {{1{{{4{b1}}}}},{{2{a2}},{a3,b5}},{1{{(p9|a4),{(b5<=b4)}}}}};
  assign y12 = (((p1?p12:p12)?{p11,p7,b3}:(p11?p0:p17))?{(p0?p17:p8),{b2},(p12?p2:p0)}:({b0}?{p11}:(p5?a2:p6)));
  assign y13 = (p14?a2:p3);
  assign y14 = (((a3!=p0)<{a1,b5,a3})||{((|b1)>(~|p0))});
  assign y15 = {4{{1{(-4'sd5)}}}};
  assign y16 = {{1{((&(~&(p2>=p14)))?({b0}?{4{b5}}:(&p9)):{3{(p5?p9:a2)}})}}};
  assign y17 = (-((~|(p7?p6:p9))*(p6*p11)));
endmodule
