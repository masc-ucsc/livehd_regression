module expression_00904(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{{4{(5'd8)}}}};
  localparam [4:0] p1 = ((((5'd14)*(5'sd12))^((5'd27)+(4'd6)))&((5'd2 * (4'd2))>=((-5'sd12)>>>(3'd1))));
  localparam [5:0] p2 = ((!{(5'd8),(-5'sd10)})?(3'sd1):((2'd2)^(-2'sd0)));
  localparam signed [3:0] p3 = (((2'd1)?(-4'sd3):(3'd4))?((2'sd1)>>(2'd1)):((5'sd10)<<<(3'sd3)));
  localparam signed [4:0] p4 = (&(3'sd1));
  localparam signed [5:0] p5 = {4{(-4'sd7)}};
  localparam [3:0] p6 = (((2'sd1)?(4'sd5):(5'd31))?((3'd3)?(-4'sd2):(-5'sd9)):((3'd7)?(4'd4):(-4'sd1)));
  localparam [4:0] p7 = (|(2'sd1));
  localparam [5:0] p8 = (&((|((4'd4)?(4'd13):(2'd2)))?(|(|((2'sd0)?(-3'sd1):(4'sd2)))):(~|((4'sd7)?(3'sd1):(3'd7)))));
  localparam signed [3:0] p9 = (((4'd2)?(-5'sd13):(4'sd1))?((2'd2)?(4'sd6):(3'd5)):(~|(-4'sd1)));
  localparam signed [4:0] p10 = {2{(+({3{(3'd6)}}|(^(-2'sd1))))}};
  localparam signed [5:0] p11 = ((-3'sd1)>>(2'd1));
  localparam [3:0] p12 = {3{(-2'sd0)}};
  localparam [4:0] p13 = (!(~&(-2'sd0)));
  localparam [5:0] p14 = (-4'sd7);
  localparam signed [3:0] p15 = (((5'd20)<(3'd1))<<<(!(-4'sd4)));
  localparam signed [4:0] p16 = (((4'd11)<<<(2'd3))?(~|(5'd3)):((3'sd3)!==(-2'sd0)));
  localparam signed [5:0] p17 = (((5'sd1)?(4'd12):(5'd24))?((2'd0)?(5'd12):(5'sd15)):{4{(2'sd1)}});

  assign y0 = {(~^(~|{(b1>>a0),(+b2),(~&b2)})),{1{((!(+a4))+(b1<b4))}},(~^({3{a5}}^~{4{b1}}))};
  assign y1 = $signed(((b5?p10:p14)?((a3?p8:b2)):(p6?p13:a2)));
  assign y2 = ((p17&p1)?(b5>>>b0):{b3,a5});
  assign y3 = ((5'd2)|$unsigned(b2));
  assign y4 = (((a2?b1:a5)?{1{b4}}:(a0<<b1))?{(b2&a4),(a1?b0:b0),(+a4)}:(-({a4,a5,b2}!={a4,a5})));
  assign y5 = ({(b2?p7:p8),(b0?p16:p4),(4'sd2)});
  assign y6 = (3'sd2);
  assign y7 = ((&(~^(~|(a1*b5))))-(^$unsigned((&(a2&&b5)))));
  assign y8 = ($unsigned(((-(~^(~&$signed((~|(~^(+$signed((^(-$unsigned($unsigned((!$signed(p9)))))))))))))))));
  assign y9 = ((|(a4>=p13))?(-(a3&&a3)):(b2?p11:p3));
  assign y10 = ({3{{{1{(4'd8)}}}}});
  assign y11 = ({((b2?a2:a5)>>>(b2))}?((a4?b0:a0)?$signed(b0):(a3>>a1)):{(b1!=a4),(a1?a0:b5),{a4,b4,a1}});
  assign y12 = ((3'sd3)^((b1!==b2)+(p2<=p15)));
  assign y13 = (|(-3'sd1));
  assign y14 = {3{(^(~|{(b5!=a3),(-a5)}))}};
  assign y15 = {(p12?p3:a3),((p15|b2)<<<(b0===a2))};
  assign y16 = (+(((a3>>b4)===(~&b5))==(&(&(p8&&b0)))));
  assign y17 = (^((b3<<p9)>(p2-a4)));
endmodule
