module expression_00291(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {(3'd2)};
  localparam [4:0] p1 = {{3{(2'sd0)}},{4{(-2'sd1)}},{4{(4'd11)}}};
  localparam [5:0] p2 = ((((2'd1)?(3'd5):(2'sd1))>>>(2'sd0))?(-2'sd1):(((4'd2)^(5'sd11))*((3'd3)!==(5'd12))));
  localparam signed [3:0] p3 = ({(((3'd1)>>(4'sd2))&((5'd9)<<<(-2'sd1)))}>>>{((-3'sd3)^~(5'd14)),{(5'd11)}});
  localparam signed [4:0] p4 = (5'd2 * (5'd12));
  localparam signed [5:0] p5 = ({{3{(2'd3)}}}||((-5'sd7)!==((2'd2)>>>(4'sd2))));
  localparam [3:0] p6 = (|(((-2'sd0)/(-5'sd7))?((3'sd3)?(2'sd0):(4'sd0)):(!(3'd4))));
  localparam [4:0] p7 = ((3'sd2)||{4{((4'sd7)>=(-5'sd11))}});
  localparam [5:0] p8 = (~|(~|{(-3'sd2),(2'd1),(3'sd3)}));
  localparam signed [3:0] p9 = {((-2'sd0)?(4'd11):(2'd2)),(^(~|(5'd16))),(2'd0)};
  localparam signed [4:0] p10 = (|(^((^((&(-3'sd3))?((3'd3)-(-3'sd0)):{2{(5'sd11)}}))^~(^({(-5'sd2)}?(^(-5'sd6)):{(5'd23)})))));
  localparam signed [5:0] p11 = (!(~|(~^(|(~&(~&(~(~|(^(~&(-2'sd1)))))))))));
  localparam [3:0] p12 = {2{{4{(5'sd9)}}}};
  localparam [4:0] p13 = (+(|(-({(|((3'sd2)<(3'd3)))}<{((2'sd1)||(3'd3)),(^(5'sd2))}))));
  localparam [5:0] p14 = ((((-2'sd1)*(4'd0))&((4'sd3)^~(3'd5)))<<((6'd2 * (2'd3))+((-3'sd1)>>>(3'sd2))));
  localparam signed [3:0] p15 = (({(4'sd5),(3'sd0)}+((2'd0)>=(2'sd0)))&&({(-2'sd1),(5'd17)}?((-2'sd0)===(3'sd1)):((5'd29)>>(3'sd1))));
  localparam signed [4:0] p16 = (~&(4'd12));
  localparam signed [5:0] p17 = (-3'sd0);

  assign y0 = (p11<=b1);
  assign y1 = (6'd2 * b1);
  assign y2 = ((!(^(~&((p0<p14)<=(p15>>>a0)))))<<<((~|{3{p15}})&((~|p17)|{p3,p8,p12})));
  assign y3 = (b2<<a4);
  assign y4 = (~^((&((p11<=a5)>(p7&&b4)))?((p3<<p10)?(p5+p13):{p6,a1,p3}):((b0?p0:p10)>(p5?p10:p1))));
  assign y5 = {(5'd23),(3'sd2)};
  assign y6 = (4'd15);
  assign y7 = ((-5'sd2)<<<(4'd2 * (2'd0)));
  assign y8 = (+{{1{({3{b4}}!=={(!(5'sd15))})}},(({a2}>>(p3?p3:b2))^~(4'sd6))});
  assign y9 = (((a0?p6:p12)?(a4<=p6):$unsigned(a1))?($signed((a4?b4:b4))||(p17-b4)):((p9?a1:b0)?(a2^p2):(p8)));
  assign y10 = (b4==p5);
  assign y11 = (((b0?b4:b4)^~{2{(b0?a3:a1)}})===(((a5<<a2))&&((a0>>>b4)&(a4&a2))));
  assign y12 = (!(~(&{3{((a1===b3)&&(a3>>a1))}})));
  assign y13 = (&(5'sd7));
  assign y14 = ((b2)&&(p5<<b1));
  assign y15 = {3{(p12>=b1)}};
  assign y16 = $unsigned($unsigned(((&$signed((b5?p10:b3)))?(-((b0^b0)<<(~&b2))):$unsigned($unsigned((a4<<<a5))))));
  assign y17 = (-4'sd2);
endmodule
