module expression_00344(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((2'd3)?(5'sd10):(2'd0));
  localparam [4:0] p1 = {4{(2'd3)}};
  localparam [5:0] p2 = (((4'd4)&(5'sd2))-(2'd3));
  localparam signed [3:0] p3 = {1{(((3'd6)<(2'd0))>=((4'd3)+(2'd0)))}};
  localparam signed [4:0] p4 = ((((-5'sd15)?(-2'sd0):(5'sd2))?((4'sd7)&&(5'd31)):((-3'sd0)!==(-5'sd9)))|(((-3'sd1)?(-4'sd0):(3'sd1))||((4'sd3)?(-5'sd6):(5'd14))));
  localparam signed [5:0] p5 = ((-4'sd1)<(2'sd0));
  localparam [3:0] p6 = (^((2'd1)?(4'd14):(5'd23)));
  localparam [4:0] p7 = {2{({4{(-4'sd0)}}^((2'd3)>>(-3'sd0)))}};
  localparam [5:0] p8 = (((~&{(2'sd0),(2'd1)})^~{((5'd24)^~(2'd0)),(&(2'd3))})|{(+((5'd2 * (3'd2))||(~^(|(-5'sd6)))))});
  localparam signed [3:0] p9 = {4{(-5'sd4)}};
  localparam signed [4:0] p10 = (|(~((-2'sd1)===(3'd2))));
  localparam signed [5:0] p11 = ((((5'd1)?(-5'sd12):(5'sd7))>>>{4{(-2'sd1)}})?((2'd2)?(-3'sd0):(-4'sd2)):((3'd7)?(-4'sd4):(2'sd0)));
  localparam [3:0] p12 = ((2'sd1)||(-2'sd1));
  localparam [4:0] p13 = (4'd2 * ((2'd3)!=(3'd7)));
  localparam [5:0] p14 = {2{(4'sd2)}};
  localparam signed [3:0] p15 = (4'd2);
  localparam signed [4:0] p16 = {3{(-2'sd1)}};
  localparam signed [5:0] p17 = {{1{{1{((3'sd2)&&(-5'sd5))}}}},{4{(2'd3)}},({(2'd3),(-5'sd3),(-3'sd1)}+((2'd2)>=(2'd2)))};

  assign y0 = (-3'sd2);
  assign y1 = (!(p16>>>b3));
  assign y2 = (-2'sd1);
  assign y3 = ({(~^a5)}?(~&(|b5)):(a4?b3:a3));
  assign y4 = {a0};
  assign y5 = ((5'd17)+(~^{3{b2}}));
  assign y6 = {p12,b1};
  assign y7 = (((p7<b2)<<(p3+p9))||((p14||p6)|{(p2|p16)}));
  assign y8 = (3'sd0);
  assign y9 = ((a3?a3:b4)!==({1{b2}}===(a2<<a3)));
  assign y10 = {2{(~^(~&((p3?p8:b4)?{3{p6}}:(a2?p5:p10))))}};
  assign y11 = (-4'sd0);
  assign y12 = ({1{({4{p17}}<<<(p12<=p6))}}?((p7?p0:p1)<<(p7^~p11)):{2{(p16?p6:p8)}});
  assign y13 = ($signed({{a4,a4,b3},(b2?b1:b0)})?$signed({(b2?a4:a2)}):((a3?b2:a0)));
  assign y14 = (!((^((~b2)>=(~|b5)))>=((b1^~b2)!=(~(b0>b5)))));
  assign y15 = ((p11?p11:p6)<(+(~^p12)));
  assign y16 = (a1?a0:b0);
  assign y17 = ((b5>>p12)?(-(^p2)):(~^(b2?b3:b2)));
endmodule
