module expression_00250(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((^((-2'sd1)===(5'sd2)))<<((2'd3)>>(-4'sd6)));
  localparam [4:0] p1 = (((2'sd0)?(3'sd1):(3'd2))?((-3'sd0)?(3'd7):(-5'sd1)):((4'sd0)?(-4'sd3):(4'sd7)));
  localparam [5:0] p2 = (^(((5'sd13)&&(3'd1))>>>(&(-4'sd2))));
  localparam signed [3:0] p3 = (!{({(2'd0),(5'sd3)}>{(3'd6),(2'd2)}),({(2'sd1),(-3'sd0)}>>{(2'd2),(3'd4),(2'd2)})});
  localparam signed [4:0] p4 = ((-(((5'd1)?(2'd2):(-2'sd1))<((4'd2)?(5'd25):(5'sd1))))-(~|(~^((5'd28)===(4'd2)))));
  localparam signed [5:0] p5 = {(&(|(~((3'sd3)?(5'd14):(3'd2))))),({(3'sd0),(3'd4)}?((-5'sd3)?(4'd2):(2'd3)):{(-2'sd1)}),(((3'd4)?(5'd16):(-2'sd1))?{(4'd2)}:((4'd15)?(2'd2):(3'sd2)))};
  localparam [3:0] p6 = ({(4'd7),(2'd3),(3'sd3)}>>>{1{{(-4'sd0),(3'd7),(3'd1)}}});
  localparam [4:0] p7 = {1{((-3'sd3)?{4{(3'd2)}}:{4{(-5'sd13)}})}};
  localparam [5:0] p8 = (((2'd2)?(-3'sd2):(2'd1))?((3'sd0)?(-5'sd14):(4'd1)):((2'sd1)?(2'sd1):(4'd1)));
  localparam signed [3:0] p9 = {{(((3'd4)+(3'sd1))+((5'd27)<<(3'sd2))),({4{(2'd0)}}^~{(4'sd0),(2'd1)})}};
  localparam signed [4:0] p10 = (!{2{{2{((5'd6)?(3'sd3):(2'd0))}}}});
  localparam signed [5:0] p11 = ((((4'd12)?(2'd0):(5'd23))?{3{(-2'sd1)}}:{4{(4'd8)}})!==(6'd2 * ((2'd2)?(4'd7):(5'd3))));
  localparam [3:0] p12 = ((!(-((-4'sd3)<<<(2'd0))))?(!((2'sd1)-(2'sd0))):((3'sd1)?(-3'sd0):(-3'sd1)));
  localparam [4:0] p13 = ((5'sd6)?(3'sd3):(-3'sd0));
  localparam [5:0] p14 = ((((4'sd6)?(4'sd1):(3'd1))/(2'sd1))^((5'd2 * (4'd13))&&(^((2'd1)?(-2'sd1):(5'd17)))));
  localparam signed [3:0] p15 = (2'sd0);
  localparam signed [4:0] p16 = ((((5'd29)?(4'd2):(2'd3))?(~^(4'd1)):((2'sd0)?(4'sd7):(5'd12)))===(((3'd0)>>(2'd2))&((-4'sd5)<<<(4'd15))));
  localparam signed [5:0] p17 = {1{{2{{3{(5'd4)}}}}}};

  assign y0 = ((~^(&p8))*(~|$unsigned(p9)));
  assign y1 = ((p12?p1:p16)/p2);
  assign y2 = {3{({2{a2}}!==(+b0))}};
  assign y3 = (!((6'd2 * (~(+a2)))>>>((b0<<<p0)+(b4<<<p13))));
  assign y4 = {1{({2{(p3||a4)}}^{(b0+b3),(-a3),(~|b0)})}};
  assign y5 = ((~^((a5?p8:a1)?(b5?a3:p4):(a2|p7)))>>((a3||a2)===(b3?a1:b4)));
  assign y6 = {(p15?p10:p12),((p3==p10)^{p9,p17,p2}),{(p16?p6:p10)}};
  assign y7 = (~((~&$signed(b4))===(^(a5|a3))));
  assign y8 = (+((a5<=b0)?(&p11):(p13?p3:p17)));
  assign y9 = (~^(4'd5));
  assign y10 = {{1{(~&(&p3))}},((p4?p14:p2)<{p5}),(&(+{2{p10}}))};
  assign y11 = (((p17?p1:b4)?(!b5):(p7&a1))^((p1<b3)==(a0&b5)));
  assign y12 = (-((5'd2 * $unsigned((a0<p0)))>=(((p16/a4))-(a0*a1))));
  assign y13 = (^{$signed((({a4,a0}!=(b1<b2))!==(+(b5===a2))))});
  assign y14 = $signed((~&(3'd5)));
  assign y15 = (4'd2 * (5'd2 * a2));
  assign y16 = (4'd2 * {3{p8}});
  assign y17 = (-(b5==p10));
endmodule
