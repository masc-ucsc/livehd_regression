module expression_00868(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{4{(4'd2)}},{1{(~|(-5'sd13))}}};
  localparam [4:0] p1 = {2{(~|((2'd2)+(3'sd0)))}};
  localparam [5:0] p2 = (&{3{(-(4'd12))}});
  localparam signed [3:0] p3 = {((-(-5'sd1))-(~|(4'sd2))),(|(|(~(&(5'd2))))),(~^{((4'sd1)&(4'd8))})};
  localparam signed [4:0] p4 = (~^(~^(3'sd0)));
  localparam signed [5:0] p5 = ({((3'd6)-(4'sd7)),((5'd9)==(5'sd11))}>>(((-5'sd7)>>(2'd2))>>>{(|(4'sd3))}));
  localparam [3:0] p6 = {4{{(4'd3),(5'sd10),(4'd10)}}};
  localparam [4:0] p7 = (~(|(((~(3'd3))>=(~&(3'd6)))<((~|(-3'sd3))==((2'sd0)&(4'sd2))))));
  localparam [5:0] p8 = (((5'sd6)?(3'sd1):(4'sd4))&&(&(4'd15)));
  localparam signed [3:0] p9 = (({1{(2'd0)}}<((-3'sd1)<(5'd14)))>>>(!(~&(((3'd2)^(5'sd14))>>((-4'sd5)?(-3'sd3):(4'sd1))))));
  localparam signed [4:0] p10 = {4{(5'sd6)}};
  localparam signed [5:0] p11 = (((5'd26)>(5'd0))*((3'd3)||(2'sd1)));
  localparam [3:0] p12 = ({4{(3'd0)}}?{4{(2'd3)}}:{4{(3'd1)}});
  localparam [4:0] p13 = (+(~&{((~&(4'd0))?(|(2'd2)):(~(3'sd0))),(-{(~^(4'sd1)),(|(3'd4)),((-5'sd9)?(3'd3):(5'd7))})}));
  localparam [5:0] p14 = (~|(!(&(~|(-(+(~(3'd7))))))));
  localparam signed [3:0] p15 = ((((3'sd1)||(-4'sd6))===(5'sd9))^(-5'sd0));
  localparam signed [4:0] p16 = (((4'd3)?(4'd9):(3'sd1))<<<((5'sd14)?(-3'sd1):(3'd6)));
  localparam signed [5:0] p17 = (~&((((5'sd3)?(2'd0):(-5'sd2))?((4'd0)?(-3'sd0):(3'd5)):(&(-2'sd1)))===((+(-2'sd0))>=((-2'sd1)<<<(-3'sd2)))));

  assign y0 = (2'd2);
  assign y1 = (5'd10);
  assign y2 = ((4'd3));
  assign y3 = {{((p13)>={4{p10}}),((a2>=b2)!=={b4,a2,b4})},{3{{b3,a0}}}};
  assign y4 = {(b2?a5:b5)};
  assign y5 = {3{(b4&&a4)}};
  assign y6 = {3{{4{p14}}}};
  assign y7 = ((~&((a4>=b1)^(a0&&b3)))!==((5'd2 * a1)&&(~&(b1==a2))));
  assign y8 = ((3'sd1)>>(($signed(p11))));
  assign y9 = ((a5*b3)^~$signed(p6));
  assign y10 = ({{p17,p10,p7},(p3?p16:p13)}?{3{p15}}:(p6?p10:p10));
  assign y11 = ((+p12)?(-3'sd0):(+p17));
  assign y12 = (6'd2 * (4'd11));
  assign y13 = (({3{b5}}?(a4?b2:b4):(5'sd0))^((a5?p15:b3)^(b1?a1:a2)));
  assign y14 = (((a3==b5)+(5'd17))&&{(b4&a0),(b4+b5),(b3?b1:a2)});
  assign y15 = (((5'd21)|{p12,p11})>>(((5'd11))&&{3{p11}}));
  assign y16 = (~($signed((3'd3))/p6));
  assign y17 = ($signed({3{$signed($unsigned(p6))}}));
endmodule
