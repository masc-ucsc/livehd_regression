module expression_00944(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (~&{4{((2'sd0)===(2'sd0))}});
  localparam [4:0] p1 = ((((3'd1)>(2'd3))?((2'sd0)!==(3'd2)):((5'd28)?(4'd1):(2'd1)))>>(2'sd0));
  localparam [5:0] p2 = ((((3'd3)?(5'sd13):(4'd10))+((3'd4)?(2'd3):(2'd3)))>(+(~(^{{{4{(4'd14)}}}}))));
  localparam signed [3:0] p3 = ((-4'sd1)<<(5'd21));
  localparam signed [4:0] p4 = ((4'd8)&(5'd24));
  localparam signed [5:0] p5 = (|(-{4{(^(~|(5'd11)))}}));
  localparam [3:0] p6 = (!(-(2'd1)));
  localparam [4:0] p7 = ({3{((4'd4)?(-5'sd6):(2'sd0))}}?(!{1{{1{{1{(3'd0)}}}}}}):(4'sd3));
  localparam [5:0] p8 = (+(((3'd5)?(-4'sd5):(5'd0))?((5'd1)<<(2'd0)):((-3'sd0)&&(-3'sd1))));
  localparam signed [3:0] p9 = (2'd3);
  localparam signed [4:0] p10 = (5'd17);
  localparam signed [5:0] p11 = ((((2'd2)&(3'sd3))<(2'd3))<<(((5'sd3)+(2'd2))!={(2'sd0),(-2'sd0),(5'd31)}));
  localparam [3:0] p12 = {2{(-2'sd0)}};
  localparam [4:0] p13 = (((3'sd1)?(4'd13):(2'sd0))?(3'd4):((-4'sd4)?(5'd18):(4'sd3)));
  localparam [5:0] p14 = (((!(3'd1))&(~(3'd3)))<<(-((4'd12)-(4'sd3))));
  localparam signed [3:0] p15 = (^(5'sd5));
  localparam signed [4:0] p16 = (|{(~|{(!(3'd2))}),(~&(!(^(4'sd4))))});
  localparam signed [5:0] p17 = {3{(^((2'd3)-(2'd0)))}};

  assign y0 = (~^p16);
  assign y1 = (^{(((^p6)^~(p11&a2))^(4'd14))});
  assign y2 = ((((a0?b3:b0)>>>{4{b2}})!=={1{{4{b3}}}})&&{2{{3{(a3?p5:a3)}}}});
  assign y3 = ($signed((3'd7))&(((2'sd0)^(p6))>>((a2<=b5)<<<(p13>=p14))));
  assign y4 = ({(p17||a3)}>=($unsigned((b1))));
  assign y5 = (({3{p14}}?$unsigned(p17):(p12>>>p13))==({2{p13}}&&(p8>=p13)));
  assign y6 = (((~&(6'd2 * b1))===(!(^(~&b0))))|(^{{{b0,b2,a3},{b1,b3,p5},(&a4)}}));
  assign y7 = ({b1,a3}!==(a2?b1:b5));
  assign y8 = (^p3);
  assign y9 = (a0?b2:b0);
  assign y10 = ((b1?b1:b3)?(p14?b1:b5):(b3?b5:a4));
  assign y11 = ((!b5)&&(p10&p6));
  assign y12 = {2{p5}};
  assign y13 = (~&(-{(~&(~^(~^(p1?p12:p3)))),{$unsigned((^{p13}))}}));
  assign y14 = ((a3==a0)?{3{a3}}:{3{b2}});
  assign y15 = ({(~{p5}),{p17,p16}}?(+(~|(-{{p4},{p9,p1}}))):{(p5?p8:p3),(+p16),(&p7)});
  assign y16 = {$unsigned(((a4?p13:p10)>>{a2,a5})),(-((4'sd5)?$unsigned(p8):(~&b3)))};
  assign y17 = ((((4'sd2)>=(p0+p1))<((+b4)|(3'd3)))&(((a5>=a2)&(p8>p1))||((p10==p15)<(-5'sd3))));
endmodule
