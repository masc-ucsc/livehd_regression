module expression_00571(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {2{(((4'd6)>=(5'd31))-((3'd7)<(2'd3)))}};
  localparam [4:0] p1 = (^((((-5'sd15)!==(4'd10))||((2'sd0)==(2'd1)))^((4'd2 * (5'd19))<(~((-2'sd1)<<<(3'd2))))));
  localparam [5:0] p2 = (&({3{{3{(5'd25)}}}}&(((5'd17)+(4'sd6))==(|{(3'd5),(2'sd0)}))));
  localparam signed [3:0] p3 = ((((-2'sd0)^(3'd5))-{(3'sd0),(5'd10),(4'd14)})^(((2'd1)>>(-5'sd12))&((3'sd1)<=(5'd24))));
  localparam signed [4:0] p4 = (!((4'sd3)^(-2'sd1)));
  localparam signed [5:0] p5 = ((((5'd3)?(3'sd3):(4'd11))?{(5'd21),(2'd3)}:{(5'd23),(5'd30),(5'sd1)})<(((5'd13)&&(5'd0))<((2'sd1)?(3'd7):(5'd2))));
  localparam [3:0] p6 = (4'd8);
  localparam [4:0] p7 = {{{{{(-5'sd7)}},((-3'sd0)!==(5'd10))},{{((4'd7)>>(2'sd0))},((4'sd7)>>>(-4'sd7))}}};
  localparam [5:0] p8 = (({1{(3'd6)}}&((3'sd0)?(-2'sd1):(5'd31)))!==(5'd9));
  localparam signed [3:0] p9 = (({3{(3'd5)}}?(~(4'sd4)):(+(5'sd10)))>=((~{4{(-4'sd4)}})^(~((5'sd7)?(2'd3):(-5'sd10)))));
  localparam signed [4:0] p10 = {4{({4{(2'd3)}}>={4{(5'd20)}})}};
  localparam signed [5:0] p11 = ((((2'd1)^(5'd3))<<((3'sd2)<<(3'd7)))>{((-2'sd1)-(-3'sd3))});
  localparam [3:0] p12 = {{{{{(2'd0),(5'sd14),(2'sd1)}},(~|(~^(5'sd0))),{(3'sd2),(2'd3)}}}};
  localparam [4:0] p13 = (!((~^(~{(4'd9),(4'sd5),(3'sd1)}))^{(+{(5'sd9),(-5'sd12),(-4'sd2)})}));
  localparam [5:0] p14 = (5'd10);
  localparam signed [3:0] p15 = (&((~|((&(~&(3'sd1)))*(^(|(2'sd1)))))===((~&((-4'sd6)&&(4'sd0)))<((5'd25)-(-5'sd2)))));
  localparam signed [4:0] p16 = ((-3'sd3)%(4'sd6));
  localparam signed [5:0] p17 = (2'd0);

  assign y0 = ($unsigned(p12)^~$unsigned(p9));
  assign y1 = (2'd1);
  assign y2 = $signed(p1);
  assign y3 = (~^(&(-4'sd3)));
  assign y4 = ((+(^(~b1)))?(b1?b4:p8):(p17?b2:a2));
  assign y5 = (b3==a0);
  assign y6 = (b4&b2);
  assign y7 = (p9>>>p7);
  assign y8 = (~&(|(&(-3'sd2))));
  assign y9 = ((b4==p7)&(p12<b0));
  assign y10 = (+((-5'sd0)?(2'd1):$unsigned(p15)));
  assign y11 = ((&(2'd3))|(|((~(2'd0))!==((5'd29)))));
  assign y12 = {(b4?p0:p17)};
  assign y13 = ($signed((((p0>=a1)*$signed(p14))>=(~|(b0===b1))))<=((~(p2^~p17))*(5'd25)));
  assign y14 = (((a2?a2:p15)?(p10?p5:p17):(p0?p16:p14))>((b5>p11)?(p8/p15):(p17!=p9)));
  assign y15 = (((a2&&a0)&{(b2||a3)})==={((b2-a5)?{b1,b2,a4}:(b5-a0))});
  assign y16 = (~{2{{(^(!{(p16+a2)}))}}});
  assign y17 = ($unsigned((-(~|$signed({p16,p6}))))?(^{(~|p9),(p9?p6:p8),{p5,p16,p4}}):{(&{(p14?p17:p14),(^p6)})});
endmodule
