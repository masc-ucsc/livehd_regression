module expression_00682(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((-5'sd2)==(4'd2 * (2'd2)));
  localparam [4:0] p1 = (3'd5);
  localparam [5:0] p2 = ((-3'sd0)/(2'sd1));
  localparam signed [3:0] p3 = ({3{(3'd0)}}<<<(&{4{(-2'sd0)}}));
  localparam signed [4:0] p4 = {{3{(-5'sd0)}},{2{(4'd4)}}};
  localparam signed [5:0] p5 = ((2'sd1)>=(5'd28));
  localparam [3:0] p6 = (((-4'sd2)?(2'sd0):(2'sd0))>((2'sd1)?(5'd7):(3'd6)));
  localparam [4:0] p7 = ((~&(5'sd10))?(-4'sd1):(2'sd0));
  localparam [5:0] p8 = ((((3'sd0)%(5'd18))?((4'd11)%(-3'sd2)):(~|(2'd0)))>((4'd4)?(~^(3'sd2)):((2'd2)!==(4'd11))));
  localparam signed [3:0] p9 = ({3{{1{(4'd7)}}}}|(~&(^((2'sd0)?(-4'sd1):(2'd3)))));
  localparam signed [4:0] p10 = {{4{{(-5'sd7)}}},{1{(((4'sd6)>=(-5'sd0))?{(3'd5)}:((5'sd4)?(2'd1):(-5'sd2)))}}};
  localparam signed [5:0] p11 = {{4{((-2'sd0)^(-2'sd1))}}};
  localparam [3:0] p12 = ({((5'sd1)||(-5'sd8))}<<<{{2{(5'sd15)}}});
  localparam [4:0] p13 = (((5'd14)?(3'sd3):(5'd29))-{1{((4'd6)<=(2'd0))}});
  localparam [5:0] p14 = (((2'd0)?(3'd6):{(5'd20)})|{((4'sd6)||(3'sd3)),((5'd0)&&(2'd3))});
  localparam signed [3:0] p15 = (-(+((5'd30)>>>(4'sd4))));
  localparam signed [4:0] p16 = {3{(-5'sd4)}};
  localparam signed [5:0] p17 = (~|(~(~^(~{(^{(4'd12),(2'd2)}),(~&(2'sd1))}))));

  assign y0 = ((((p0<<a3)-({p17,b5}))^((a5+a1)>>(5'd2 * b0))));
  assign y1 = (~(~((p0<<<a0)*(a5&&a4))));
  assign y2 = {((~&(a5!=p17))<(p2|a5)),(~{{p14,p11},(|a3)}),((p6!=a3)|{b5,p2})};
  assign y3 = (5'sd5);
  assign y4 = (-(^$unsigned((+(!(~^$signed($signed(((^(~(~&a2))))))))))));
  assign y5 = ((p16?b0:b5)?(b3&p7):(b5>>>b3));
  assign y6 = (a0!==a2);
  assign y7 = ({1{(b0?p17:a4)}}?(p1>=p9):(p5^a0));
  assign y8 = (((b1>=b4)==(a1/b3))>=((b1)<<<(a2&&b0)));
  assign y9 = ((!(|$signed(((a2<p15)>=(~^b2)))))|(&(~|(~|(~^(b3===b3))))));
  assign y10 = {1{(~(!(-3'sd2)))}};
  assign y11 = (-(({b0,b4,a4})===$signed((|{(b2<<<a2)}))));
  assign y12 = {1{{3{b0}}}};
  assign y13 = ((+(b3?a0:p7))<$unsigned((~^(p8))));
  assign y14 = (~^{a2,b1,b0});
  assign y15 = ((!(~|((p13)^~(~&b4))))||((~|(a0||b2))%a1));
  assign y16 = (-((p16<p2)?(b3===b2):(4'd2 * p14)));
  assign y17 = {p7,p13,p2};
endmodule
