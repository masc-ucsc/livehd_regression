module expression_00613(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (-{2{{4{(2'd2)}}}});
  localparam [4:0] p1 = (3'sd3);
  localparam [5:0] p2 = {{3{(3'd0)}},(-2'sd0)};
  localparam signed [3:0] p3 = {(4'd6),(5'd20),(2'sd1)};
  localparam signed [4:0] p4 = (~^((-2'sd1)^~(-4'sd0)));
  localparam signed [5:0] p5 = ((~&(((-5'sd4)+(2'sd0))+((4'd7)+(4'd13))))>=(6'd2 * ((5'd15)>>(2'd1))));
  localparam [3:0] p6 = (((3'd0)^~(4'd13))>>>((2'd3)^(5'sd15)));
  localparam [4:0] p7 = {2{{4{(2'd1)}}}};
  localparam [5:0] p8 = (((5'd28)|(5'sd4))?((-2'sd0)?(4'd1):(3'd0)):((-4'sd2)|(5'd8)));
  localparam signed [3:0] p9 = (((-4'sd6)<<<(5'd11))>(((-5'sd5)+(2'd3))*(-((-2'sd0)!=(-5'sd13)))));
  localparam signed [4:0] p10 = {2{(5'd24)}};
  localparam signed [5:0] p11 = ((&((3'sd0)!=(3'd7)))|((2'd1)?(-2'sd0):(3'd5)));
  localparam [3:0] p12 = (-5'sd11);
  localparam [4:0] p13 = {(({1{(3'd6)}}||{(2'd3)})>>({(4'd7),(2'sd0),(3'd0)}<<<{(5'sd8),(5'd29)}))};
  localparam [5:0] p14 = ((((3'sd2)||(4'd14))===((3'd1)||(4'sd1)))===((-3'sd1)>>(+(-5'sd7))));
  localparam signed [3:0] p15 = {{(2'd0)}};
  localparam signed [4:0] p16 = ({4{(2'd1)}}^(|(3'sd3)));
  localparam signed [5:0] p17 = {2{(4'sd4)}};

  assign y0 = (~|((-4'sd1)>(3'sd1)));
  assign y1 = {3{{2{(a4||p13)}}}};
  assign y2 = {4{({2{b4}}^(-2'sd0))}};
  assign y3 = ({2{((5'sd11))}}!=(5'd2 * {4{b2}}));
  assign y4 = (4'sd2);
  assign y5 = $unsigned(b0);
  assign y6 = ((+((b5<b2)===(a1&a5)))<((p5&&p4)>>>(b3<<p13)));
  assign y7 = (-3'sd3);
  assign y8 = ({3{{p12,p4}}}<=(~^(5'd0)));
  assign y9 = (($unsigned((+(a1<<<a3)))==((a4==p2)^(5'sd11)))^~({2{(&a4)}}||((|b5)<=(b1!==b3))));
  assign y10 = (|(-4'sd6));
  assign y11 = (((p14)*(a4))<<<$unsigned((|(~|(~^p10)))));
  assign y12 = (((!(&p6))<<(a0===a2))+{{3{a1}},{2{p13}},(p8^a0)});
  assign y13 = ({{p2,p10,p12}}||(|(~&{p13,p15,a0})));
  assign y14 = (~|(-3'sd1));
  assign y15 = $unsigned($unsigned((~&$unsigned((4'd11)))));
  assign y16 = (&((!((4'd2 * $unsigned((~a4)))))<=(~&((-(~(a0<a0)))<<<$unsigned($unsigned((~|a1)))))));
  assign y17 = {((~^p6)+(p16==a1)),(~(~&(p11-p5))),{b5,a2,p4}};
endmodule
