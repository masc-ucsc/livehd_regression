module expression_00382(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = (((2'sd0)?(3'd3):(4'd3))<=((3'sd0)<<<(4'sd2)));
  localparam [4:0] p1 = (~{1{((2'd0)==(-4'sd5))}});
  localparam [5:0] p2 = (((-5'sd10)>=(4'd0))^~{(3'd4),(5'd31),(3'd5)});
  localparam signed [3:0] p3 = (&{4{{2{(-3'sd3)}}}});
  localparam signed [4:0] p4 = ((5'd4)<<(5'd0));
  localparam signed [5:0] p5 = (((5'd3)==(-2'sd0))^~((-5'sd10)-(-4'sd0)));
  localparam [3:0] p6 = {4{((2'd0)?(-5'sd14):(4'd4))}};
  localparam [4:0] p7 = ({((3'sd2)?(2'd3):(-4'sd4)),(!(4'sd5)),((-2'sd0)?(2'd1):(2'd0))}>(~{1{(~&((2'sd1)?(-5'sd14):(2'd0)))}}));
  localparam [5:0] p8 = {{{(^(2'd2)),{(3'd2),(5'sd13)}},(~^(!(+(3'sd1))))},(~^(^{(~^(!{{(-3'sd0),(4'd5),(2'd1)}}))}))};
  localparam signed [3:0] p9 = ((5'd20)&(((5'sd8)+(2'sd1))?((2'sd0)/(5'sd6)):(2'sd1)));
  localparam signed [4:0] p10 = (((2'd3)+(2'sd0))>>>(-3'sd0));
  localparam signed [5:0] p11 = (!({1{((-2'sd0)?(-4'sd1):(5'sd11))}}>{1{((-5'sd0)?(5'd25):(2'd2))}}));
  localparam [3:0] p12 = (+((!(4'd2 * (5'd22)))===((4'd13)-(2'd3))));
  localparam [4:0] p13 = {3{(3'd6)}};
  localparam [5:0] p14 = (((5'sd11)%(3'd0))&((4'd2)==(4'd7)));
  localparam signed [3:0] p15 = ((-2'sd1)?{(-5'sd1),(3'sd0)}:(5'd31));
  localparam signed [4:0] p16 = (((3'sd3)?(4'd11):(5'd24))?(5'd2 * ((5'd0)<=(3'd0))):{3{(-4'sd7)}});
  localparam signed [5:0] p17 = (~^({(2'sd1),(4'sd4)}+((3'd2)^~(3'sd3))));

  assign y0 = (~&{(p14<p2),(p5<p1)});
  assign y1 = ((a0?p14:a4)?(p8?b0:a4):(a3<<<p1));
  assign y2 = ((b1?b2:b5)?(~a4):(&p14));
  assign y3 = ({{a5,p13},(p7>=b5),(b5<<a2)}^{4{a0}});
  assign y4 = (!({4{a3}}-(p12&b2)));
  assign y5 = {4{{1{{4{b3}}}}}};
  assign y6 = $signed((^{4{(&(p8>>p4))}}));
  assign y7 = (+(({1{p16}}<<<(p12<<p2))&&((p12|p7)&&(!p16))));
  assign y8 = (~^({1{(p7-p7)}}<=((p1!=p5)<=(p3<p12))));
  assign y9 = {1{(~|((b1===a4)?(3'd2):(^(p15<<<b0))))}};
  assign y10 = ((6'd2 * (b1<=p12))^~((p6>=p1)*(p11-p9)));
  assign y11 = (((p17>>a1)>>(3'd0))?({p13}?(a1===b2):(~|p4)):{{(4'd13),(a4==p13)}});
  assign y12 = $unsigned((((((&b0))&&{{2{b2}}})||{{2{b2}},(a5>=b2),(a4!=p2)})));
  assign y13 = {{{$signed(((a4?a1:p2)|(&p3)))}},$signed(((b5?p16:a5)||(~&(p1?a1:p8))))};
  assign y14 = {{3{$unsigned(p16)}},$signed(((b2+p16)?{2{b3}}:(b0===a3))),(4'sd0)};
  assign y15 = (-(~^{1{({3{a0}}>=(b3?p17:a3))}}));
  assign y16 = (~|a3);
  assign y17 = ({4{b3}}?(a2?p3:p12):{4{p4}});
endmodule
