module expression_00896(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((5'd2 * (2'd0))>(5'd16));
  localparam [4:0] p1 = (~|((6'd2 * ((5'd3)<<<(2'd3)))>(6'd2 * ((5'd1)|(5'd27)))));
  localparam [5:0] p2 = (-(-{4{(+{2{(5'd23)}})}}));
  localparam signed [3:0] p3 = (({(4'd10),(3'sd2),(5'd2)}+(-(3'd7)))<=(!(-{(2'd0),(-4'sd3)})));
  localparam signed [4:0] p4 = (&((-((-5'sd8)?(3'sd2):(4'd10)))?(-((-4'sd7)*(2'd3))):(^((5'sd9)>>>(4'd6)))));
  localparam signed [5:0] p5 = {2{(3'd6)}};
  localparam [3:0] p6 = ({{(4'sd7),(4'd11),(-2'sd0)},(3'd2),{(5'sd15)}}-({2{(-3'sd1)}}^~(-2'sd0)));
  localparam [4:0] p7 = (2'sd0);
  localparam [5:0] p8 = (&(~^(-((((4'd9)!==(2'sd0))>(4'd10))+{4{(3'sd3)}}))));
  localparam signed [3:0] p9 = {2{{(~|(-2'sd1))}}};
  localparam signed [4:0] p10 = {4{(!((2'd0)&&(5'sd5)))}};
  localparam signed [5:0] p11 = {1{(+{4{{1{((3'd5)==(3'd7))}}}})}};
  localparam [3:0] p12 = {3{((4'd9)?(-3'sd2):(3'd1))}};
  localparam [4:0] p13 = ((((4'd2)!=(4'd4))?((5'sd0)>=(-4'sd1)):((3'd4)+(-4'sd5)))^~(((-5'sd3)&(4'd1))===((-3'sd1)!=(2'd0))));
  localparam [5:0] p14 = (({1{(2'd0)}}?((-3'sd1)>=(3'sd1)):((4'd2)<<(5'd11)))^~(((4'd1)!==(5'sd5))!=((5'd15)?(4'd5):(3'd3))));
  localparam signed [3:0] p15 = (((+(~^(3'sd3)))^((5'sd3)!==(4'd2)))<<((~&(^(-5'sd4)))<(~|(-(-4'sd4)))));
  localparam signed [4:0] p16 = {2{{2{(5'sd1)}}}};
  localparam signed [5:0] p17 = {(!(~|(4'sd1)))};

  assign y0 = (~|(~&{1{{4{b1}}}}));
  assign y1 = (^$unsigned((^$signed({4{(-b3)}}))));
  assign y2 = ($unsigned(((5'sd1)&&(6'd2 * a0)))<=($unsigned(b3)==(~|b1)));
  assign y3 = {(~|(!{{(-p3),(^p3)}}))};
  assign y4 = {1{$signed((~^($signed(((p6<p13)?(p1?p4:b5):(p9?p4:p1)))>=(({2{p6}}^~{3{p10}})))))}};
  assign y5 = ({3{(b4===b5)}}!==(-(~((a2^b2)>=(a2>=a4)))));
  assign y6 = ((5'sd8)?$signed((p3?p12:p16)):((+p0)|(p6<<p15)));
  assign y7 = (~^(((a0>>>p10)?(a3?b5:b0):(~a3))+(|(~^(5'd29)))));
  assign y8 = {(!{p7,p7,b5}),(p15^a4),{(~|p9)}};
  assign y9 = (5'd2 * (~^(p12<p0)));
  assign y10 = {(((a4&&b5)=={1{b3}})-((p14<<a3)-{b5}))};
  assign y11 = ((-($unsigned(p6)/b3))<=((+a4)+(p15%p2)));
  assign y12 = {3{(~^{1{{2{$signed(p9)}}}})}};
  assign y13 = {2{b1}};
  assign y14 = {((p3?p12:p13)?{p2,p9,a2}:(p13?p4:p15))};
  assign y15 = {{{{p6,p14,p12},(p1?p10:p5),(p3<p17)},{2{(p15?p0:p12)}}}};
  assign y16 = {(-$signed(((p14)))),(~(~^(|(p5?p5:p1))))};
  assign y17 = ({1{(a2!=b2)}}&&{4{p9}});
endmodule
