module expression_00158(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {3{((4'd13)|(-5'sd2))}};
  localparam [4:0] p1 = (~|{{(-2'sd1),(-2'sd0)},{(3'sd2),(2'd2),(3'd7)},{(-2'sd0),(-5'sd14)}});
  localparam [5:0] p2 = ((3'd1)>=((^((2'sd1)^(-2'sd1)))>>(5'd12)));
  localparam signed [3:0] p3 = {2{{2{(-3'sd0)}}}};
  localparam signed [4:0] p4 = ((((5'sd2)>>>(2'd1))^~(&(-(5'sd10))))^(-4'sd5));
  localparam signed [5:0] p5 = (((5'd7)>=(-2'sd1))?((3'd3)?(4'd3):(2'sd0)):((5'd21)?(4'd0):(-2'sd0)));
  localparam [3:0] p6 = (~|((5'sd15)?(-5'sd6):(2'd2)));
  localparam [4:0] p7 = {{4{{(5'sd11),(3'd6),(5'sd12)}}},(|(2'd2))};
  localparam [5:0] p8 = ((-4'sd3)<<(-2'sd1));
  localparam signed [3:0] p9 = ((3'd2)&(-4'sd1));
  localparam signed [4:0] p10 = (~|{((5'sd3)?(-3'sd3):(3'sd1))});
  localparam signed [5:0] p11 = ((2'd0)<<(3'd6));
  localparam [3:0] p12 = ((5'd13)>>(5'sd2));
  localparam [4:0] p13 = {((-4'sd4)&&{(3'sd0)}),(~|{(-(4'sd7))})};
  localparam [5:0] p14 = (^({(3'd4),(5'sd15),(2'd3)}!=={(+(3'd3)),(!(3'd3))}));
  localparam signed [3:0] p15 = ((-(+((-2'sd1)|(-2'sd0))))&&(((4'sd1)>(-2'sd1))<=((5'd28)==(5'd5))));
  localparam signed [4:0] p16 = ((2'd3)>(3'sd0));
  localparam signed [5:0] p17 = (((4'd1)>=(3'sd3))?(3'd3):((3'd4)==(4'sd0)));

  assign y0 = (({3{a5}}?(p13>>>b1):{1{p15}})?({{p2,p11}}>{4{p14}}):({2{b3}}?(4'd2 * b0):(a3^~a4)));
  assign y1 = ((|{1{(5'sd10)}})^(~|(|{1{{(|(b1||p3)),(a4>p2)}}})));
  assign y2 = (^{1{(~|(((b1==a5)?(~&b2):(~a5))?{3{(~|b3)}}:{4{a5}}))}});
  assign y3 = ((&(-(~$signed((~^$signed(a0))))))>>>(-((a0+b4)||(~&(|b2)))));
  assign y4 = ($unsigned(({b2,a4,a4}?(p12?a1:a3):(a3?b0:a3)))+{($signed($unsigned((((b2?b3:a5)||(b4?b4:b0))))))});
  assign y5 = {3{(p4?p0:a5)}};
  assign y6 = (+(-(5'd27)));
  assign y7 = (+(((p12<=p15)<<(-5'sd1))^(+(3'sd2))));
  assign y8 = ((a4-b2)/p4);
  assign y9 = (&({p11,p4,p1}+(~^p10)));
  assign y10 = ((^($unsigned((~&(^($unsigned(p9)))))-(~^((a3)===$unsigned(b3))))));
  assign y11 = $signed(p5);
  assign y12 = {p10,p17};
  assign y13 = {3{(~&{(~^p5),(p8&&p6),(b4>=p8)})}};
  assign y14 = ((p13?p16:a0)*(&$signed(b1)));
  assign y15 = (~|{2{(~|{2{(+{3{a5}})}})}});
  assign y16 = (({2{p4}}?(~p13):{4{p2}})?(~|((~p2)?{3{p13}}:(p9?p13:p12))):(!((p5-p6)^(p17?p13:p8))));
  assign y17 = (a1?a2:a0);
endmodule
