module expression_00370(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = {{((4'sd5)<<<(2'd1)),{(2'd3),(-4'sd7),(4'd12)},((5'd22)&(2'd3))}};
  localparam [4:0] p1 = {{4{(2'd1)}},(-(-4'sd6)),(4'd5)};
  localparam [5:0] p2 = (4'sd4);
  localparam signed [3:0] p3 = {({(2'd1),(4'sd3),(5'sd4)}?((2'sd0)?(4'd5):(3'd5)):{(3'd5)}),{((2'd3)<(4'd5)),((4'sd3)?(2'd2):(2'sd1)),{(3'sd0),(3'd2),(-4'sd2)}}};
  localparam signed [4:0] p4 = (4'd10);
  localparam signed [5:0] p5 = ((((5'd8)>(5'sd13))?(|(5'sd6)):(~|(3'd7)))?(((-2'sd1)<(4'sd7))>>((-2'sd0)/(-5'sd3))):(((-3'sd1)?(4'sd3):(4'd3))<((4'd3)||(4'd12))));
  localparam [3:0] p6 = ((((4'sd0)>>(5'sd3))<<<((5'd7)!=(3'd2)))^~(((4'd10)^~(4'd8))|((4'sd2)<<(3'sd0))));
  localparam [4:0] p7 = {4{{3{(-3'sd3)}}}};
  localparam [5:0] p8 = (3'd6);
  localparam signed [3:0] p9 = {4{(2'd2)}};
  localparam signed [4:0] p10 = ((-4'sd5)?{(3'sd1),(4'd9),(4'd4)}:((2'd2)?(3'd1):(4'd1)));
  localparam signed [5:0] p11 = (~^((!(^{(~&{(5'd8),(3'd3)})}))&&((!((5'sd4)<(-4'sd4)))||(!(|(-2'sd0))))));
  localparam [3:0] p12 = {(((2'd2)&(4'sd6))&(2'd1)),({4{(-5'sd4)}}<<{2{(2'd1)}}),(4'sd6)};
  localparam [4:0] p13 = (((&(~&(!(5'd7))))===(((4'd12)<<(4'd6))<=((3'sd1)|(4'd11))))>>>(|({1{{3{(-5'sd4)}}}}<<<{3{(-4'sd0)}})));
  localparam [5:0] p14 = ((((3'sd1)||(4'd11))>((-3'sd0)&&(4'd8)))&((4'd6)?(5'd14):(3'sd1)));
  localparam signed [3:0] p15 = {3{({2{(4'd8)}}|((5'd25)^(2'sd1)))}};
  localparam signed [4:0] p16 = (~^(~(^(&(2'd2)))));
  localparam signed [5:0] p17 = (~|(3'sd3));

  assign y0 = (2'd2);
  assign y1 = (-((~^$signed($signed(((b2<<<p6)?(^b1):(a4)))))||(^(~$signed((-(b2?a3:b2)))))));
  assign y2 = (!{(~^(!(5'd2 * $unsigned($signed(p3)))))});
  assign y3 = {1{(~|(3'd2))}};
  assign y4 = {3{(~^$unsigned((~&(6'd2 * b1))))}};
  assign y5 = {({(5'd15)}+{p14,b5,a3}),((^(p8<<<p8))||({a4,b5}===(2'd2)))};
  assign y6 = ({4{p17}}|(5'sd9));
  assign y7 = {1{(p15<=p0)}};
  assign y8 = (2'sd1);
  assign y9 = {2{p0}};
  assign y10 = ((4'd1)-((p15<<<p10)<$unsigned((4'd13))));
  assign y11 = ((~p8)<{4{p1}});
  assign y12 = {2{{1{((~^b2)<(p10?b1:p2))}}}};
  assign y13 = {4{{1{(b5^~p4)}}}};
  assign y14 = (&{3{(!(+(b5-b1)))}});
  assign y15 = (4'd12);
  assign y16 = {4{(p2^a5)}};
  assign y17 = {{(~(~|b3))},{a1,b5,a5},(^(&(!a2)))};
endmodule
