module expression_00577(a0, a1, a2, a3, a4, a5, b0, b1, b2, b3, b4, b5, y);
  input [3:0] a0;
  input [4:0] a1;
  input [5:0] a2;
  input signed [3:0] a3;
  input signed [4:0] a4;
  input signed [5:0] a5;

  input [3:0] b0;
  input [4:0] b1;
  input [5:0] b2;
  input signed [3:0] b3;
  input signed [4:0] b4;
  input signed [5:0] b5;

  wire [3:0] y0;
  wire [4:0] y1;
  wire [5:0] y2;
  wire signed [3:0] y3;
  wire signed [4:0] y4;
  wire signed [5:0] y5;
  wire [3:0] y6;
  wire [4:0] y7;
  wire [5:0] y8;
  wire signed [3:0] y9;
  wire signed [4:0] y10;
  wire signed [5:0] y11;
  wire [3:0] y12;
  wire [4:0] y13;
  wire [5:0] y14;
  wire signed [3:0] y15;
  wire signed [4:0] y16;
  wire signed [5:0] y17;

  output [89:0] y;
  assign y = {y0,y1,y2,y3,y4,y5,y6,y7,y8,y9,y10,y11,y12,y13,y14,y15,y16,y17};

  localparam [3:0] p0 = ((~(5'd23))>>>(~^(3'd0)));
  localparam [4:0] p1 = (~{3{((-2'sd0)<=(3'd0))}});
  localparam [5:0] p2 = (4'd2 * ((3'd7)<<(4'd14)));
  localparam signed [3:0] p3 = ((|({3{(4'd0)}}=={2{(2'd1)}}))-(~^(-{2{{1{(2'd0)}}}})));
  localparam signed [4:0] p4 = ((4'd9)^(-4'sd4));
  localparam signed [5:0] p5 = (({{(-3'sd1),(5'd25)}}^((3'sd3)&&(5'd18)))&&(((4'sd7)>(3'd0))-((2'sd1)||(4'd14))));
  localparam [3:0] p6 = (~^((((5'd7)>>(4'sd2))>>>((3'sd1)?(-2'sd0):(2'sd0)))^~(^(~^(((5'd18)?(2'sd1):(5'd26))&&((-2'sd0)?(2'd2):(4'sd0)))))));
  localparam [4:0] p7 = (~|(((3'd1)?(-5'sd10):(2'd2))*((4'sd6)>(3'sd2))));
  localparam [5:0] p8 = (((((2'sd1)&(3'd0))&&((5'sd13)>>>(5'd5)))&&(((5'd5)%(4'd15))&&((-5'sd13)<<<(4'sd3))))<(((5'd13)>(3'd0))/(-2'sd1)));
  localparam signed [3:0] p9 = ({((-4'sd1)&(3'd6))}|(~&(^(-4'sd7))));
  localparam signed [4:0] p10 = ((-2'sd1)?(3'sd0):(3'sd0));
  localparam signed [5:0] p11 = {1{{((2'sd0)?(2'sd0):(-2'sd0)),((-2'sd1)>>>(2'd0)),((-5'sd3)>=(-2'sd1))}}};
  localparam [3:0] p12 = {(-3'sd0),(2'd1)};
  localparam [4:0] p13 = (~^((((3'sd3)!==(2'd0))|((-5'sd3)>>>(2'd1)))&({4{(-3'sd0)}}+((5'd19)-(3'sd3)))));
  localparam [5:0] p14 = (+(3'sd0));
  localparam signed [3:0] p15 = ((4'd2 * (!((2'd1)?(2'd3):(3'd6))))==(({(4'd8)}&((4'd11)?(3'd6):(3'd2)))-(~^((-4'sd2)?(5'sd1):(4'd4)))));
  localparam signed [4:0] p16 = (5'd11);
  localparam signed [5:0] p17 = ({3{(2'd1)}}?(~&{(2'd2),(-5'sd1)}):(2'd2));

  assign y0 = (|((~(+(-(~(b1?a0:b1)))))?((~|p9)?(-p11):(|p15)):((p11?a1:a0)?(~p5):(+b3))));
  assign y1 = (~^({(a0?a1:b0),(4'd13),{a4}}==={(-4'sd5),(b1!=a1)}));
  assign y2 = (!(^{($signed((b3||a0))?(5'd2 * b0):(a1>=a4)),((~{b1})?(a5<<<a0):(p7<<a0))}));
  assign y3 = (-5'sd6);
  assign y4 = (a2?a1:p12);
  assign y5 = (!$signed((!{({p10,b2}>(6'd2 * a0)),({p0,b4,a5}|(~^(a3>=a4)))})));
  assign y6 = (p7&p7);
  assign y7 = ((-2'sd0));
  assign y8 = ((!(4'sd4))-((b1?b0:b2)?(&b4):(&b5)));
  assign y9 = ((-{2{(~^{1{(^a4)}})}})<<<{4{(+b2)}});
  assign y10 = (4'd5);
  assign y11 = ($unsigned((2'sd1))?$unsigned(((a3?a3:b1))):(~(&(&(5'd0)))));
  assign y12 = (3'd5);
  assign y13 = (((a0&&b4)||(p3&a4))<<<((b5<a0)|(p12>>>p8)));
  assign y14 = {(2'd1),(p16?p11:a0)};
  assign y15 = (((((b3)||(b3<=a5)))+$signed({(p11>b4)}))<<(((a3==a5)<(a1!==b4))!==$signed(({b0}<<(b3+b0)))));
  assign y16 = (((2'd0)<(p7?p16:p0))+$signed((p5?p14:b0)));
  assign y17 = ({(p6?p0:b1),(a0?p3:p9)}>(~(^(a1==p4))));
endmodule
